version https://git-lfs.github.com/spec/v1
oid sha256:99c02a2898ecdd52de5c9a4a7461b10445ea25d436b1645b2a20574a1f4dd966
size 344049
