# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2014, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *       NGLibraryCreator, Development_version_64 - build 201405300513        *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on us19.nangate.us for user Lucio Rech (lre).
# Local time is now Tue, 3 Jun 2014, 13:07:07.
# Main process id is 12480.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2_X1_8T
  CLASS core ;
  FOREIGN AND2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.4639 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0847 0.078 0.35 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.076 0.334 0.4267 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.108 0.1419 0.1267 ;
        RECT 0.114 0.1267 0.1419 0.2853 ;
        RECT 0.114 0.2853 0.1419 0.3627 ;
        RECT 0.1419 0.108 0.242 0.1267 ;
        RECT 0.242 0.108 0.27 0.1267 ;
        RECT 0.242 0.1267 0.27 0.2853 ;
      LAYER M1 ;
        RECT 0.114 0.108 0.1419 0.1267 ;
        RECT 0.114 0.1267 0.1419 0.2853 ;
        RECT 0.114 0.2853 0.1419 0.3627 ;
        RECT 0.1419 0.108 0.242 0.1267 ;
        RECT 0.242 0.108 0.27 0.1267 ;
        RECT 0.242 0.1267 0.27 0.2853 ;
  END
END AND2_X1_8T

MACRO AND2_X2_8T
  CLASS core ;
  FOREIGN AND2_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.1653 0.083 0.3467 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.0427 0.306 0.0867 ;
        RECT 0.302 0.4253 0.306 0.4693 ;
        RECT 0.306 0.0427 0.334 0.0867 ;
        RECT 0.306 0.0867 0.334 0.4253 ;
        RECT 0.306 0.4253 0.334 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.3827 0.082 0.4013 ;
        RECT 0.082 0.1107 0.242 0.1293 ;
        RECT 0.082 0.3827 0.242 0.4013 ;
        RECT 0.242 0.1107 0.27 0.1293 ;
        RECT 0.242 0.1293 0.27 0.3827 ;
        RECT 0.242 0.3827 0.27 0.4013 ;
      LAYER M1 ;
        RECT 0.054 0.3827 0.082 0.4013 ;
        RECT 0.082 0.1107 0.242 0.1293 ;
        RECT 0.082 0.3827 0.242 0.4013 ;
        RECT 0.242 0.1107 0.27 0.1293 ;
        RECT 0.242 0.1293 0.27 0.3827 ;
        RECT 0.242 0.3827 0.27 0.4013 ;
  END
END AND2_X2_8T

MACRO AND3_X1_8T
  CLASS core ;
  FOREIGN AND3_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.128 0.334 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1729 0.128 0.211 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.128 0.08 0.384 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.076 0.462 0.436 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.079 0.0667 0.238 0.066732 ;
        RECT 0.054 0.4207 0.274 0.4393 ;
        RECT 0.274 0.0633 0.37 0.0913 ;
        RECT 0.274 0.4207 0.37 0.4393 ;
        RECT 0.37 0.0633 0.398 0.0913 ;
        RECT 0.37 0.0913 0.398 0.4207 ;
        RECT 0.37 0.4207 0.398 0.4393 ;
      LAYER M1 ;
        RECT 0.079 0.0667 0.238 0.066732 ;
        RECT 0.054 0.4207 0.274 0.4393 ;
        RECT 0.274 0.0633 0.37 0.0913 ;
        RECT 0.274 0.4207 0.37 0.4393 ;
        RECT 0.37 0.0633 0.398 0.0913 ;
        RECT 0.37 0.0913 0.398 0.4207 ;
        RECT 0.37 0.4207 0.398 0.4393 ;
  END
END AND3_X1_8T

MACRO AND3_X2_8T
  CLASS core ;
  FOREIGN AND3_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.2133 0.206 0.342 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.1707 0.083 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2013 0.27 0.358 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.366 0.0427 0.37 0.1047 ;
        RECT 0.366 0.4253 0.37 0.4693 ;
        RECT 0.37 0.0427 0.398 0.1047 ;
        RECT 0.37 0.1047 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.048 0.08 0.104 ;
        RECT 0.048 0.104 0.08 0.1253 ;
        RECT 0.08 0.104 0.298 0.1253 ;
        RECT 0.054 0.3873 0.146 0.4087 ;
        RECT 0.146 0.1493 0.306 0.168 ;
        RECT 0.146 0.3873 0.306 0.4087 ;
        RECT 0.306 0.1493 0.334 0.168 ;
        RECT 0.306 0.168 0.334 0.3873 ;
        RECT 0.306 0.3873 0.334 0.4087 ;
      LAYER M1 ;
        RECT 0.048 0.048 0.08 0.104 ;
        RECT 0.048 0.104 0.08 0.1253 ;
        RECT 0.08 0.104 0.298 0.1253 ;
        RECT 0.054 0.3873 0.146 0.4087 ;
        RECT 0.146 0.1493 0.306 0.168 ;
        RECT 0.146 0.3873 0.306 0.4087 ;
        RECT 0.306 0.1493 0.334 0.168 ;
        RECT 0.306 0.168 0.334 0.3873 ;
        RECT 0.306 0.3873 0.334 0.4087 ;
  END
END AND3_X2_8T

MACRO AND4_X1_8T
  CLASS core ;
  FOREIGN AND4_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.128 0.398 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.128 0.272 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.128 0.1419 0.3413 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.076 0.526 0.436 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.462 0.5307 ;
        RECT 0.462 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.424 0.338 0.4453 ;
        RECT 0.338 0.0667 0.434 0.066732 ;
        RECT 0.338 0.424 0.434 0.4453 ;
        RECT 0.434 0.0667 0.462 0.066732 ;
        RECT 0.434 0.088 0.462 0.424 ;
        RECT 0.434 0.424 0.462 0.4453 ;
        RECT 0.1409 0.066 0.298 0.098 ;
      LAYER M1 ;
        RECT 0.082 0.424 0.338 0.4453 ;
        RECT 0.338 0.0667 0.434 0.066732 ;
        RECT 0.338 0.424 0.434 0.4453 ;
        RECT 0.434 0.0667 0.462 0.066732 ;
        RECT 0.434 0.088 0.462 0.424 ;
        RECT 0.434 0.424 0.462 0.4453 ;
        RECT 0.1409 0.066 0.298 0.098 ;
  END
END AND4_X1_8T

MACRO AND4_X2_8T
  CLASS core ;
  FOREIGN AND4_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.1607 0.398 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.128 0.27 0.3847 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.128 0.1419 0.3847 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.3847 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.064 0.526 0.4267 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.462 0.5307 ;
        RECT 0.462 0.4933 0.65 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.65 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0667419 0.0667 0.298 0.066732 ;
        RECT 0.082 0.424 0.342 0.4453 ;
        RECT 0.342 0.11 0.434 0.1313 ;
        RECT 0.342 0.424 0.434 0.4453 ;
        RECT 0.434 0.11 0.462 0.1313 ;
        RECT 0.434 0.1313 0.462 0.424 ;
        RECT 0.434 0.424 0.462 0.4453 ;
      LAYER M1 ;
        RECT 0.0667419 0.0667 0.298 0.066732 ;
        RECT 0.082 0.424 0.342 0.4453 ;
        RECT 0.342 0.11 0.434 0.1313 ;
        RECT 0.342 0.424 0.434 0.4453 ;
        RECT 0.434 0.11 0.462 0.1313 ;
        RECT 0.434 0.1313 0.462 0.424 ;
        RECT 0.434 0.424 0.462 0.4453 ;
  END
END AND4_X2_8T

MACRO ANTENNA_8T
  CLASS core ;
  FOREIGN ANTENNA_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
END ANTENNA_8T

MACRO AOI21_X1_8T
  CLASS core ;
  FOREIGN AOI21_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.128 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0893 0.078 0.3413 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.128 0.334 0.3413 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.066714 0.0667 0.0667419 0.066732 ;
        RECT 0.114 0.088 0.1419 0.3573 ;
        RECT 0.0667419 0.0667 0.306 0.066732 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.298 0.5307 ;
        RECT 0.298 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.3867 0.08 0.408 ;
        RECT 0.048 0.408 0.08 0.4693 ;
        RECT 0.08 0.3867 0.298 0.408 ;
      LAYER M1 ;
        RECT 0.048 0.3867 0.08 0.408 ;
        RECT 0.048 0.408 0.08 0.4693 ;
        RECT 0.08 0.3867 0.298 0.408 ;
  END
END AOI21_X1_8T

MACRO AOI21_X2_8T
  CLASS core ;
  FOREIGN AOI21_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.2013 0.398 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1533 0.27 0.172 ;
        RECT 0.242 0.172 0.27 0.2987 ;
        RECT 0.242 0.2987 0.27 0.3413 ;
        RECT 0.27 0.1533 0.493 0.172 ;
        RECT 0.493 0.1533 0.531 0.172 ;
        RECT 0.493 0.172 0.531 0.2987 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.2987 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.077 0.1107 0.178 0.1293 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.326 ;
        RECT 0.178 0.326 0.206 0.3806 ;
        RECT 0.178 0.3806 0.206 0.3993 ;
        RECT 0.206 0.1107 0.43 0.1293 ;
        RECT 0.206 0.3806 0.43 0.3993 ;
        RECT 0.43 0.3806 0.434 0.3993 ;
        RECT 0.434 0.326 0.462 0.3806 ;
        RECT 0.434 0.3806 0.462 0.3993 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.535 0.5307 ;
        RECT 0.535 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.3667 0.08 0.4233 ;
        RECT 0.048 0.4233 0.08 0.446 ;
        RECT 0.08 0.4233 0.498 0.446 ;
        RECT 0.498 0.344 0.526 0.3667 ;
        RECT 0.498 0.3667 0.526 0.4233 ;
        RECT 0.498 0.4233 0.526 0.446 ;
        RECT 0.146 0.0679 0.535 0.0867 ;
      LAYER M1 ;
        RECT 0.048 0.3667 0.08 0.4233 ;
        RECT 0.048 0.4233 0.08 0.446 ;
        RECT 0.08 0.4233 0.498 0.446 ;
        RECT 0.498 0.344 0.526 0.3667 ;
        RECT 0.498 0.3667 0.526 0.4233 ;
        RECT 0.498 0.4233 0.526 0.446 ;
        RECT 0.146 0.0679 0.535 0.0867 ;
  END
END AOI21_X2_8T

MACRO AOI22_X1_8T
  CLASS core ;
  FOREIGN AOI22_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.128 0.27 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.128 0.398 0.3233 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.132 0.1419 0.384 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1409 0.0679 0.306 0.0867 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.0867 0.334 0.388 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.42 0.37 0.4493 ;
        RECT 0.37 0.3687 0.398 0.42 ;
        RECT 0.37 0.42 0.398 0.4493 ;
      LAYER M1 ;
        RECT 0.082 0.42 0.37 0.4493 ;
        RECT 0.37 0.3687 0.398 0.42 ;
        RECT 0.37 0.42 0.398 0.4493 ;
  END
END AOI22_X1_8T

MACRO AOI22_X2_8T
  CLASS core ;
  FOREIGN AOI22_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.1827 0.462 0.2013 ;
        RECT 0.434 0.2013 0.462 0.326 ;
        RECT 0.434 0.326 0.462 0.3413 ;
        RECT 0.462 0.1827 0.654 0.2013 ;
        RECT 0.654 0.1827 0.6899 0.2013 ;
        RECT 0.6899 0.1827 0.718 0.2013 ;
        RECT 0.6899 0.2013 0.718 0.326 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.2467 0.59 0.3413 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.204 0.204 0.334 0.3507 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1613 0.078 0.3413 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.133342 0.1333 0.13337 0.133328 ;
        RECT 0.242 0.152 0.27 0.1527 ;
        RECT 0.242 0.1527 0.27 0.2133 ;
        RECT 0.13337 0.1333 0.362 0.133328 ;
        RECT 0.362 0.1333 0.37 0.133328 ;
        RECT 0.37 0.1333 0.398 0.133328 ;
        RECT 0.37 0.152 0.398 0.1527 ;
        RECT 0.37 0.1527 0.398 0.2133 ;
        RECT 0.37 0.2133 0.398 0.3087 ;
        RECT 0.37 0.3087 0.398 0.3786 ;
        RECT 0.37 0.3786 0.398 0.4013 ;
        RECT 0.398 0.1333 0.626 0.133328 ;
        RECT 0.398 0.152 0.626 0.1527 ;
        RECT 0.398 0.3786 0.626 0.4013 ;
        RECT 0.626 0.1333 0.654 0.133328 ;
        RECT 0.626 0.152 0.654 0.1527 ;
        RECT 0.626 0.3087 0.654 0.3786 ;
        RECT 0.626 0.3786 0.654 0.4013 ;
        RECT 0.654 0.1333 0.6899 0.133328 ;
        RECT 0.654 0.152 0.6899 0.1527 ;
        RECT 0.6899 0.064 0.718 0.1333 ;
        RECT 0.6899 0.1333 0.718 0.133328 ;
        RECT 0.6899 0.152 0.718 0.1527 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.718 0.5307 ;
        RECT 0.718 0.4933 0.778 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.778 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.406 0.088 0.626 0.1093 ;
        RECT 0.626 0.048 0.654 0.088 ;
        RECT 0.626 0.088 0.654 0.1093 ;
        RECT 0.077 0.4253 0.6899 0.444 ;
        RECT 0.6899 0.3713 0.718 0.4253 ;
        RECT 0.6899 0.4253 0.718 0.444 ;
        RECT 0.0859 0.0579 0.362 0.0967 ;
      LAYER M1 ;
        RECT 0.406 0.088 0.626 0.1093 ;
        RECT 0.626 0.048 0.654 0.088 ;
        RECT 0.626 0.088 0.654 0.1093 ;
        RECT 0.077 0.4253 0.6899 0.444 ;
        RECT 0.6899 0.3713 0.718 0.4253 ;
        RECT 0.6899 0.4253 0.718 0.444 ;
        RECT 0.0859 0.0579 0.362 0.0967 ;
  END
END AOI22_X2_8T

MACRO BUF_X1_8T
  CLASS core ;
  FOREIGN BUF_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.076 0.272 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1429 0.5307 ;
        RECT 0.1429 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.048 0.115 0.1233 ;
        RECT 0.114 0.1233 0.115 0.142 ;
        RECT 0.114 0.2853 0.115 0.304 ;
        RECT 0.114 0.304 0.115 0.372 ;
        RECT 0.115 0.048 0.1419 0.1233 ;
        RECT 0.115 0.1233 0.1419 0.142 ;
        RECT 0.115 0.142 0.1419 0.2853 ;
        RECT 0.115 0.2853 0.1419 0.304 ;
        RECT 0.115 0.304 0.1419 0.372 ;
        RECT 0.1419 0.1233 0.1429 0.142 ;
        RECT 0.1419 0.142 0.1429 0.2853 ;
        RECT 0.1419 0.2853 0.1429 0.304 ;
      LAYER M1 ;
        RECT 0.114 0.048 0.115 0.1233 ;
        RECT 0.114 0.1233 0.115 0.142 ;
        RECT 0.114 0.2853 0.115 0.304 ;
        RECT 0.114 0.304 0.115 0.372 ;
        RECT 0.115 0.048 0.1419 0.1233 ;
        RECT 0.115 0.1233 0.1419 0.142 ;
        RECT 0.115 0.142 0.1419 0.2853 ;
        RECT 0.115 0.2853 0.1419 0.304 ;
        RECT 0.115 0.304 0.1419 0.372 ;
        RECT 0.1419 0.1233 0.1429 0.142 ;
        RECT 0.1419 0.142 0.1429 0.2853 ;
        RECT 0.1419 0.2853 0.1429 0.304 ;
  END
END BUF_X1_8T

MACRO BUF_X2_8T
  CLASS core ;
  FOREIGN BUF_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.178 0.078 0.3413 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1739 0.402 0.177 0.4693 ;
        RECT 0.177 0.048 0.178 0.088 ;
        RECT 0.177 0.402 0.178 0.4693 ;
        RECT 0.178 0.048 0.206 0.088 ;
        RECT 0.178 0.088 0.206 0.402 ;
        RECT 0.178 0.402 0.206 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.042 0.3707 0.05 0.3893 ;
        RECT 0.042 0.3893 0.05 0.4573 ;
        RECT 0.05 0.064 0.078 0.128 ;
        RECT 0.05 0.128 0.078 0.1467 ;
        RECT 0.05 0.3707 0.078 0.3893 ;
        RECT 0.05 0.3893 0.078 0.4573 ;
        RECT 0.078 0.128 0.0859 0.1467 ;
        RECT 0.078 0.3707 0.0859 0.3893 ;
        RECT 0.078 0.3893 0.0859 0.4573 ;
        RECT 0.0859 0.128 0.114 0.1467 ;
        RECT 0.0859 0.3707 0.114 0.3893 ;
        RECT 0.114 0.128 0.1419 0.1467 ;
        RECT 0.114 0.1467 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
      LAYER M1 ;
        RECT 0.042 0.3707 0.05 0.3893 ;
        RECT 0.042 0.3893 0.05 0.4573 ;
        RECT 0.05 0.064 0.078 0.128 ;
        RECT 0.05 0.128 0.078 0.1467 ;
        RECT 0.05 0.3707 0.078 0.3893 ;
        RECT 0.05 0.3893 0.078 0.4573 ;
        RECT 0.078 0.128 0.0859 0.1467 ;
        RECT 0.078 0.3707 0.0859 0.3893 ;
        RECT 0.078 0.3893 0.0859 0.4573 ;
        RECT 0.0859 0.128 0.114 0.1467 ;
        RECT 0.0859 0.3707 0.114 0.3893 ;
        RECT 0.114 0.128 0.1419 0.1467 ;
        RECT 0.114 0.1467 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
  END
END BUF_X2_8T

MACRO BUF_X4_8T
  CLASS core ;
  FOREIGN BUF_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1613 0.206 0.3507 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.0679 0.21 0.0867 ;
        RECT 0.21 0.0679 0.27 0.0867 ;
        RECT 0.21 0.4253 0.27 0.444 ;
        RECT 0.27 0.0679 0.368 0.0867 ;
        RECT 0.27 0.4253 0.368 0.444 ;
        RECT 0.368 0.0679 0.4 0.0867 ;
        RECT 0.368 0.0867 0.4 0.4253 ;
        RECT 0.368 0.4253 0.4 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.027 0.1107 0.0859 0.132 ;
        RECT 0.0859 0.1107 0.242 0.132 ;
        RECT 0.0859 0.3799 0.242 0.4013 ;
        RECT 0.242 0.1107 0.27 0.132 ;
        RECT 0.242 0.132 0.27 0.3799 ;
        RECT 0.242 0.3799 0.27 0.4013 ;
      LAYER M1 ;
        RECT 0.027 0.1107 0.0859 0.132 ;
        RECT 0.0859 0.1107 0.242 0.132 ;
        RECT 0.0859 0.3799 0.242 0.4013 ;
        RECT 0.242 0.1107 0.27 0.132 ;
        RECT 0.242 0.132 0.27 0.3799 ;
        RECT 0.242 0.3799 0.27 0.4013 ;
  END
END BUF_X4_8T

MACRO BUF_X8_8T
  CLASS core ;
  FOREIGN BUF_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.244 ;
        RECT 0.05 0.244 0.078 0.2653 ;
        RECT 0.05 0.2653 0.078 0.3413 ;
        RECT 0.078 0.244 0.298 0.2653 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.0679 0.7 0.0867 ;
        RECT 0.338 0.4253 0.7 0.444 ;
        RECT 0.7 0.0679 0.754 0.0867 ;
        RECT 0.7 0.4253 0.754 0.444 ;
        RECT 0.754 0.0679 0.782 0.0867 ;
        RECT 0.754 0.0867 0.782 0.4253 ;
        RECT 0.754 0.4253 0.782 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.7 0.5307 ;
        RECT 0.7 0.4933 0.906 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.906 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.099 0.0653 0.114 0.124 ;
        RECT 0.099 0.124 0.114 0.1427 ;
        RECT 0.114 0.0653 0.1419 0.124 ;
        RECT 0.114 0.124 0.1419 0.1427 ;
        RECT 0.114 0.3513 0.1419 0.3887 ;
        RECT 0.114 0.3887 0.1419 0.4467 ;
        RECT 0.1419 0.0653 0.157 0.124 ;
        RECT 0.1419 0.124 0.157 0.1427 ;
        RECT 0.1419 0.3513 0.157 0.3887 ;
        RECT 0.157 0.124 0.354 0.1427 ;
        RECT 0.157 0.3513 0.354 0.3887 ;
        RECT 0.354 0.124 0.382 0.1427 ;
        RECT 0.354 0.1427 0.382 0.2273 ;
        RECT 0.354 0.2273 0.382 0.246 ;
        RECT 0.354 0.246 0.382 0.3513 ;
        RECT 0.354 0.3513 0.382 0.3887 ;
        RECT 0.382 0.2273 0.7 0.246 ;
      LAYER M1 ;
        RECT 0.099 0.0653 0.114 0.124 ;
        RECT 0.099 0.124 0.114 0.1427 ;
        RECT 0.114 0.0653 0.1419 0.124 ;
        RECT 0.114 0.124 0.1419 0.1427 ;
        RECT 0.114 0.3513 0.1419 0.3887 ;
        RECT 0.114 0.3887 0.1419 0.4467 ;
        RECT 0.1419 0.0653 0.157 0.124 ;
        RECT 0.1419 0.124 0.157 0.1427 ;
        RECT 0.1419 0.3513 0.157 0.3887 ;
        RECT 0.157 0.124 0.354 0.1427 ;
        RECT 0.157 0.3513 0.354 0.3887 ;
        RECT 0.354 0.124 0.382 0.1427 ;
        RECT 0.354 0.1427 0.382 0.2273 ;
        RECT 0.354 0.2273 0.382 0.246 ;
        RECT 0.354 0.246 0.382 0.3513 ;
        RECT 0.354 0.3513 0.382 0.3887 ;
        RECT 0.382 0.2273 0.7 0.246 ;
  END
END BUF_X8_8T

MACRO BUF_X12_8T
  CLASS core ;
  FOREIGN BUF_X12_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.28 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.1573 0.08 0.244 ;
        RECT 0.048 0.244 0.08 0.2653 ;
        RECT 0.048 0.2653 0.08 0.3433 ;
        RECT 0.08 0.244 0.426 0.2653 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.0679 1.07 0.0867 ;
        RECT 0.466 0.4253 1.07 0.444 ;
        RECT 1.07 0.0679 1.1359 0.0867 ;
        RECT 1.07 0.4253 1.1359 0.444 ;
        RECT 1.1359 0.0679 1.168 0.0867 ;
        RECT 1.1359 0.0867 1.168 0.4253 ;
        RECT 1.1359 0.4253 1.168 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.07 0.5307 ;
        RECT 1.07 0.4933 1.29 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.29 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.098 0.3673 0.112 0.3887 ;
        RECT 0.098 0.3887 0.112 0.4467 ;
        RECT 0.112 0.0653 0.144 0.1233 ;
        RECT 0.112 0.1233 0.144 0.1447 ;
        RECT 0.112 0.3673 0.144 0.3887 ;
        RECT 0.112 0.3887 0.144 0.4467 ;
        RECT 0.144 0.1233 0.157 0.1447 ;
        RECT 0.144 0.3673 0.157 0.3887 ;
        RECT 0.144 0.3887 0.157 0.4467 ;
        RECT 0.157 0.1233 0.462 0.1447 ;
        RECT 0.157 0.3673 0.462 0.3887 ;
        RECT 0.462 0.1233 0.49 0.1447 ;
        RECT 0.462 0.1447 0.49 0.2467 ;
        RECT 0.462 0.2467 0.49 0.2653 ;
        RECT 0.462 0.2653 0.49 0.3673 ;
        RECT 0.462 0.3673 0.49 0.3887 ;
        RECT 0.49 0.2467 1.07 0.2653 ;
      LAYER M1 ;
        RECT 0.098 0.3673 0.112 0.3887 ;
        RECT 0.098 0.3887 0.112 0.4467 ;
        RECT 0.112 0.0653 0.144 0.1233 ;
        RECT 0.112 0.1233 0.144 0.1447 ;
        RECT 0.112 0.3673 0.144 0.3887 ;
        RECT 0.112 0.3887 0.144 0.4467 ;
        RECT 0.144 0.1233 0.157 0.1447 ;
        RECT 0.144 0.3673 0.157 0.3887 ;
        RECT 0.144 0.3887 0.157 0.4467 ;
        RECT 0.157 0.1233 0.462 0.1447 ;
        RECT 0.157 0.3673 0.462 0.3887 ;
        RECT 0.462 0.1233 0.49 0.1447 ;
        RECT 0.462 0.1447 0.49 0.2467 ;
        RECT 0.462 0.2467 0.49 0.2653 ;
        RECT 0.462 0.2653 0.49 0.3673 ;
        RECT 0.462 0.3673 0.49 0.3887 ;
        RECT 0.49 0.2467 1.07 0.2653 ;
  END
END BUF_X12_8T

MACRO BUF_X16_8T
  CLASS core ;
  FOREIGN BUF_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1547 0.078 0.2367 ;
        RECT 0.05 0.2367 0.078 0.2753 ;
        RECT 0.05 0.2753 0.078 0.3413 ;
        RECT 0.078 0.2367 0.554 0.2753 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.0679 1.454 0.0867 ;
        RECT 0.594 0.4213 1.454 0.44 ;
        RECT 1.454 0.0679 1.52 0.0867 ;
        RECT 1.454 0.4213 1.52 0.44 ;
        RECT 1.52 0.0679 1.552 0.0867 ;
        RECT 1.52 0.0867 1.552 0.4213 ;
        RECT 1.52 0.4213 1.552 0.44 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.454 0.5307 ;
        RECT 1.454 0.4933 1.674 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.674 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.0653 0.1419 0.1367 ;
        RECT 0.114 0.1367 0.1419 0.1553 ;
        RECT 0.114 0.3053 0.1419 0.324 ;
        RECT 0.114 0.324 0.1419 0.4287 ;
        RECT 0.1419 0.1367 0.59 0.1553 ;
        RECT 0.1419 0.3053 0.59 0.324 ;
        RECT 0.59 0.1367 0.618 0.1553 ;
        RECT 0.59 0.1553 0.618 0.2453 ;
        RECT 0.59 0.2453 0.618 0.264 ;
        RECT 0.59 0.264 0.618 0.3053 ;
        RECT 0.59 0.3053 0.618 0.324 ;
        RECT 0.618 0.2453 1.454 0.264 ;
      LAYER M1 ;
        RECT 0.114 0.0653 0.1419 0.1367 ;
        RECT 0.114 0.1367 0.1419 0.1553 ;
        RECT 0.114 0.3053 0.1419 0.324 ;
        RECT 0.114 0.324 0.1419 0.4287 ;
        RECT 0.1419 0.1367 0.59 0.1553 ;
        RECT 0.1419 0.3053 0.59 0.324 ;
        RECT 0.59 0.1367 0.618 0.1553 ;
        RECT 0.59 0.1553 0.618 0.2453 ;
        RECT 0.59 0.2453 0.618 0.264 ;
        RECT 0.59 0.264 0.618 0.3053 ;
        RECT 0.59 0.3053 0.618 0.324 ;
        RECT 0.618 0.2453 1.454 0.264 ;
  END
END BUF_X16_8T

MACRO CLKBUF_X1_8T
  CLASS core ;
  FOREIGN CLKBUF_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.076 0.272 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1429 0.5307 ;
        RECT 0.1429 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.048 0.115 0.1233 ;
        RECT 0.114 0.1233 0.115 0.142 ;
        RECT 0.114 0.262 0.115 0.3053 ;
        RECT 0.114 0.3053 0.115 0.3487 ;
        RECT 0.115 0.048 0.1419 0.1233 ;
        RECT 0.115 0.1233 0.1419 0.142 ;
        RECT 0.115 0.142 0.1419 0.262 ;
        RECT 0.115 0.262 0.1419 0.3053 ;
        RECT 0.115 0.3053 0.1419 0.3487 ;
        RECT 0.1419 0.1233 0.1429 0.142 ;
        RECT 0.1419 0.142 0.1429 0.262 ;
        RECT 0.1419 0.262 0.1429 0.3053 ;
      LAYER M1 ;
        RECT 0.114 0.048 0.115 0.1233 ;
        RECT 0.114 0.1233 0.115 0.142 ;
        RECT 0.114 0.262 0.115 0.3053 ;
        RECT 0.114 0.3053 0.115 0.3487 ;
        RECT 0.115 0.048 0.1419 0.1233 ;
        RECT 0.115 0.1233 0.1419 0.142 ;
        RECT 0.115 0.142 0.1419 0.262 ;
        RECT 0.115 0.262 0.1419 0.3053 ;
        RECT 0.115 0.3053 0.1419 0.3487 ;
        RECT 0.1419 0.1233 0.1429 0.142 ;
        RECT 0.1419 0.142 0.1429 0.262 ;
        RECT 0.1419 0.262 0.1429 0.3053 ;
  END
END CLKBUF_X1_8T

MACRO CLKBUF_X2_8T
  CLASS core ;
  FOREIGN CLKBUF_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1973 0.078 0.3413 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1739 0.4253 0.178 0.4693 ;
        RECT 0.178 0.048 0.206 0.4253 ;
        RECT 0.178 0.4253 0.206 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.086 0.08 0.128 ;
        RECT 0.048 0.128 0.08 0.1467 ;
        RECT 0.048 0.3707 0.08 0.3893 ;
        RECT 0.048 0.3893 0.08 0.4573 ;
        RECT 0.08 0.128 0.114 0.1467 ;
        RECT 0.08 0.3707 0.114 0.3893 ;
        RECT 0.114 0.128 0.1419 0.1467 ;
        RECT 0.114 0.1467 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
      LAYER M1 ;
        RECT 0.048 0.086 0.08 0.128 ;
        RECT 0.048 0.128 0.08 0.1467 ;
        RECT 0.048 0.3707 0.08 0.3893 ;
        RECT 0.048 0.3893 0.08 0.4573 ;
        RECT 0.08 0.128 0.114 0.1467 ;
        RECT 0.08 0.3707 0.114 0.3893 ;
        RECT 0.114 0.128 0.1419 0.1467 ;
        RECT 0.114 0.1467 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
  END
END CLKBUF_X2_8T

MACRO CLKBUF_X4_8T
  CLASS core ;
  FOREIGN CLKBUF_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1613 0.1419 0.3507 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.0679 0.205 0.0867 ;
        RECT 0.205 0.0679 0.206 0.0867 ;
        RECT 0.205 0.4253 0.206 0.444 ;
        RECT 0.206 0.0679 0.368 0.0867 ;
        RECT 0.206 0.4253 0.368 0.444 ;
        RECT 0.368 0.0679 0.4 0.0867 ;
        RECT 0.368 0.0867 0.4 0.4253 ;
        RECT 0.368 0.4253 0.4 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.041 0.1107 0.082 0.1293 ;
        RECT 0.082 0.1107 0.178 0.1293 ;
        RECT 0.082 0.3827 0.178 0.4013 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.3827 ;
        RECT 0.178 0.3827 0.206 0.4013 ;
      LAYER M1 ;
        RECT 0.041 0.1107 0.082 0.1293 ;
        RECT 0.082 0.1107 0.178 0.1293 ;
        RECT 0.082 0.3827 0.178 0.4013 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.3827 ;
        RECT 0.178 0.3827 0.206 0.4013 ;
  END
END CLKBUF_X4_8T

MACRO CLKBUF_X8_8T
  CLASS core ;
  FOREIGN CLKBUF_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.2187 ;
        RECT 0.05 0.2187 0.078 0.2373 ;
        RECT 0.05 0.2373 0.078 0.3413 ;
        RECT 0.078 0.1707 0.079 0.2187 ;
        RECT 0.078 0.2187 0.079 0.2373 ;
        RECT 0.079 0.2187 0.318 0.2373 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.0679 0.718 0.0867 ;
        RECT 0.338 0.4253 0.718 0.444 ;
        RECT 0.718 0.0679 0.754 0.0867 ;
        RECT 0.718 0.4253 0.754 0.444 ;
        RECT 0.754 0.0679 0.782 0.0867 ;
        RECT 0.754 0.0867 0.782 0.4253 ;
        RECT 0.754 0.4253 0.782 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.718 0.5307 ;
        RECT 0.718 0.4933 0.906 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.906 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.1107 0.114 0.1293 ;
        RECT 0.114 0.1107 0.1419 0.1293 ;
        RECT 0.114 0.3 0.1419 0.3213 ;
        RECT 0.114 0.3213 0.1419 0.3613 ;
        RECT 0.1419 0.1107 0.406 0.1293 ;
        RECT 0.1419 0.3 0.406 0.3213 ;
        RECT 0.406 0.1107 0.434 0.1293 ;
        RECT 0.406 0.1293 0.434 0.238 ;
        RECT 0.406 0.238 0.434 0.2767 ;
        RECT 0.406 0.2767 0.434 0.3 ;
        RECT 0.406 0.3 0.434 0.3213 ;
        RECT 0.434 0.238 0.718 0.2767 ;
      LAYER M1 ;
        RECT 0.05 0.1107 0.114 0.1293 ;
        RECT 0.114 0.1107 0.1419 0.1293 ;
        RECT 0.114 0.3 0.1419 0.3213 ;
        RECT 0.114 0.3213 0.1419 0.3613 ;
        RECT 0.1419 0.1107 0.406 0.1293 ;
        RECT 0.1419 0.3 0.406 0.3213 ;
        RECT 0.406 0.1107 0.434 0.1293 ;
        RECT 0.406 0.1293 0.434 0.238 ;
        RECT 0.406 0.238 0.434 0.2767 ;
        RECT 0.406 0.2767 0.434 0.3 ;
        RECT 0.406 0.3 0.434 0.3213 ;
        RECT 0.434 0.238 0.718 0.2767 ;
  END
END CLKBUF_X8_8T

MACRO CLKBUF_X12_8T
  CLASS core ;
  FOREIGN CLKBUF_X12_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.28 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.1587 0.083 0.224 ;
        RECT 0.045 0.224 0.083 0.2453 ;
        RECT 0.045 0.2453 0.083 0.3533 ;
        RECT 0.083 0.224 0.426 0.2453 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.0679 0.998 0.0867 ;
        RECT 0.466 0.4253 0.998 0.444 ;
        RECT 0.998 0.0679 1.1359 0.0867 ;
        RECT 0.998 0.4253 1.1359 0.444 ;
        RECT 1.1359 0.0679 1.168 0.0867 ;
        RECT 1.1359 0.0867 1.168 0.4253 ;
        RECT 1.1359 0.4253 1.168 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.998 0.5307 ;
        RECT 0.998 0.4933 1.29 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.29 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0429 0.1107 0.114 0.1293 ;
        RECT 0.114 0.1107 0.1419 0.1293 ;
        RECT 0.114 0.3667 0.1419 0.3853 ;
        RECT 0.114 0.3853 0.1419 0.4467 ;
        RECT 0.1419 0.1107 0.462 0.1293 ;
        RECT 0.1419 0.3667 0.462 0.3853 ;
        RECT 0.462 0.1107 0.49 0.1293 ;
        RECT 0.462 0.1293 0.49 0.2093 ;
        RECT 0.462 0.2093 0.49 0.2306 ;
        RECT 0.462 0.2306 0.49 0.3667 ;
        RECT 0.462 0.3667 0.49 0.3853 ;
        RECT 0.49 0.1107 0.494 0.1293 ;
        RECT 0.49 0.1293 0.494 0.2093 ;
        RECT 0.49 0.2093 0.494 0.2306 ;
        RECT 0.494 0.2093 0.998 0.2306 ;
      LAYER M1 ;
        RECT 0.0429 0.1107 0.114 0.1293 ;
        RECT 0.114 0.1107 0.1419 0.1293 ;
        RECT 0.114 0.3667 0.1419 0.3853 ;
        RECT 0.114 0.3853 0.1419 0.4467 ;
        RECT 0.1419 0.1107 0.462 0.1293 ;
        RECT 0.1419 0.3667 0.462 0.3853 ;
        RECT 0.462 0.1107 0.49 0.1293 ;
        RECT 0.462 0.1293 0.49 0.2093 ;
        RECT 0.462 0.2093 0.49 0.2306 ;
        RECT 0.462 0.2306 0.49 0.3667 ;
        RECT 0.462 0.3667 0.49 0.3853 ;
        RECT 0.49 0.1107 0.494 0.1293 ;
        RECT 0.49 0.1293 0.494 0.2093 ;
        RECT 0.49 0.2093 0.494 0.2306 ;
        RECT 0.494 0.2093 0.998 0.2306 ;
  END
END CLKBUF_X12_8T

MACRO CLKBUF_X16_8T
  CLASS core ;
  FOREIGN CLKBUF_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.148 0.078 0.2173 ;
        RECT 0.05 0.2173 0.078 0.2387 ;
        RECT 0.05 0.2387 0.078 0.3507 ;
        RECT 0.078 0.2173 0.554 0.2387 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.0579 1.454 0.0967 ;
        RECT 0.594 0.4153 1.454 0.454 ;
        RECT 1.454 0.0579 1.52 0.0967 ;
        RECT 1.454 0.4153 1.52 0.454 ;
        RECT 1.52 0.0579 1.552 0.0967 ;
        RECT 1.52 0.0967 1.552 0.4153 ;
        RECT 1.52 0.4153 1.552 0.454 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.454 0.5307 ;
        RECT 1.454 0.4933 1.674 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.674 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.0727 0.1419 0.1367 ;
        RECT 0.114 0.1367 0.1419 0.1553 ;
        RECT 0.114 0.35 0.1419 0.3753 ;
        RECT 0.114 0.3753 0.1419 0.4253 ;
        RECT 0.1419 0.1367 0.595 0.1553 ;
        RECT 0.1419 0.35 0.595 0.3753 ;
        RECT 0.595 0.1367 0.653 0.1553 ;
        RECT 0.595 0.1553 0.653 0.2107 ;
        RECT 0.595 0.2107 0.653 0.2293 ;
        RECT 0.595 0.2293 0.653 0.35 ;
        RECT 0.595 0.35 0.653 0.3753 ;
        RECT 0.653 0.2107 1.454 0.2293 ;
      LAYER M1 ;
        RECT 0.114 0.0727 0.1419 0.1367 ;
        RECT 0.114 0.1367 0.1419 0.1553 ;
        RECT 0.114 0.35 0.1419 0.3753 ;
        RECT 0.114 0.3753 0.1419 0.4253 ;
        RECT 0.1419 0.1367 0.595 0.1553 ;
        RECT 0.1419 0.35 0.595 0.3753 ;
        RECT 0.595 0.1367 0.653 0.1553 ;
        RECT 0.595 0.1553 0.653 0.2107 ;
        RECT 0.595 0.2107 0.653 0.2293 ;
        RECT 0.595 0.2293 0.653 0.35 ;
        RECT 0.595 0.35 0.653 0.3753 ;
        RECT 0.653 0.2107 1.454 0.2293 ;
  END
END CLKBUF_X16_8T

MACRO CLKGATETST_X1_8T
  CLASS core ;
  FOREIGN CLKGATETST_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.088 BY 0.512 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.6899 0.1587 0.718 0.3413 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.448 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.2133 0.078 0.448 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.01 0.064 1.038 0.436 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.366 0.5307 ;
        RECT 0.366 0.4933 0.91 0.5307 ;
        RECT 0.91 0.4933 0.974 0.5307 ;
        RECT 0.974 0.4933 1.098 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.098 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.21 0.268 0.686 0.2867 ;
        RECT 0.146 0.3107 0.522 0.3293 ;
        RECT 0.73 0.268 1.006 0.2867 ;
      LAYER MINT1 ;
        RECT 0.21 0.268 0.686 0.2867 ;
        RECT 0.146 0.3107 0.522 0.3293 ;
        RECT 0.73 0.268 1.006 0.2867 ;
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.238 0.0867 ;
        RECT 0.242 0.176 0.27 0.3607 ;
        RECT 0.37 0.1613 0.398 0.3347 ;
        RECT 0.462 0.248 0.494 0.34 ;
        RECT 0.626 0.1107 0.654 0.1293 ;
        RECT 0.626 0.1293 0.654 0.3707 ;
        RECT 0.626 0.3707 0.654 0.3947 ;
        RECT 0.654 0.1107 0.75 0.1293 ;
        RECT 0.654 0.3707 0.75 0.3947 ;
        RECT 0.75 0.1107 0.755 0.1293 ;
        RECT 0.754 0.1653 0.79 0.3087 ;
        RECT 0.754 0.3087 0.79 0.3347 ;
        RECT 0.79 0.3087 0.8179 0.3347 ;
        RECT 0.8179 0.3087 0.846 0.3347 ;
        RECT 0.8179 0.3347 0.846 0.3893 ;
        RECT 0.946 0.1507 0.974 0.3827 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.4187 ;
        RECT 0.178 0.4187 0.206 0.4507 ;
        RECT 0.206 0.1107 0.302 0.1293 ;
        RECT 0.206 0.4187 0.302 0.4507 ;
        RECT 0.302 0.4187 0.366 0.4507 ;
        RECT 0.306 0.2047 0.334 0.364 ;
        RECT 0.306 0.364 0.334 0.3827 ;
        RECT 0.334 0.364 0.558 0.3827 ;
        RECT 0.558 0.1227 0.59 0.2047 ;
        RECT 0.558 0.2047 0.59 0.364 ;
        RECT 0.558 0.364 0.59 0.3827 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.2227 ;
        RECT 0.462 0.0679 0.466 0.0867 ;
        RECT 0.466 0.0679 0.882 0.0867 ;
        RECT 0.466 0.4187 0.882 0.4507 ;
        RECT 0.882 0.0679 0.91 0.0867 ;
        RECT 0.882 0.0867 0.91 0.2227 ;
        RECT 0.882 0.2227 0.91 0.4187 ;
        RECT 0.882 0.4187 0.91 0.4507 ;
      LAYER V1 ;
        RECT 0.178 0.3107 0.206 0.3293 ;
        RECT 0.242 0.268 0.27 0.2867 ;
        RECT 0.37 0.268 0.398 0.2867 ;
        RECT 0.462 0.3107 0.49 0.3293 ;
        RECT 0.626 0.268 0.654 0.2867 ;
        RECT 0.762 0.268 0.79 0.2867 ;
        RECT 0.946 0.268 0.974 0.2867 ;
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.238 0.0867 ;
        RECT 0.242 0.176 0.27 0.3607 ;
        RECT 0.37 0.1613 0.398 0.3347 ;
        RECT 0.462 0.248 0.494 0.34 ;
        RECT 0.626 0.1107 0.654 0.1293 ;
        RECT 0.626 0.1293 0.654 0.3707 ;
        RECT 0.626 0.3707 0.654 0.3947 ;
        RECT 0.654 0.1107 0.75 0.1293 ;
        RECT 0.654 0.3707 0.75 0.3947 ;
        RECT 0.75 0.1107 0.755 0.1293 ;
        RECT 0.754 0.1653 0.79 0.3087 ;
        RECT 0.754 0.3087 0.79 0.3347 ;
        RECT 0.79 0.3087 0.8179 0.3347 ;
        RECT 0.8179 0.3087 0.846 0.3347 ;
        RECT 0.8179 0.3347 0.846 0.3893 ;
        RECT 0.946 0.1507 0.974 0.3827 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.4187 ;
        RECT 0.178 0.4187 0.206 0.4507 ;
        RECT 0.206 0.1107 0.302 0.1293 ;
        RECT 0.206 0.4187 0.302 0.4507 ;
        RECT 0.302 0.4187 0.366 0.4507 ;
        RECT 0.306 0.2047 0.334 0.364 ;
        RECT 0.306 0.364 0.334 0.3827 ;
        RECT 0.334 0.364 0.558 0.3827 ;
        RECT 0.558 0.1227 0.59 0.2047 ;
        RECT 0.558 0.2047 0.59 0.364 ;
        RECT 0.558 0.364 0.59 0.3827 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.2227 ;
        RECT 0.462 0.0679 0.466 0.0867 ;
        RECT 0.466 0.0679 0.882 0.0867 ;
        RECT 0.466 0.4187 0.882 0.4507 ;
        RECT 0.882 0.0679 0.91 0.0867 ;
        RECT 0.882 0.0867 0.91 0.2227 ;
        RECT 0.882 0.2227 0.91 0.4187 ;
        RECT 0.882 0.4187 0.91 0.4507 ;
  END
END CLKGATETST_X1_8T

MACRO DFFRNQ_X1_8T
  CLASS core ;
  FOREIGN DFFRNQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.3507 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.704 0.1827 1.1339 0.2013 ;
        RECT 1.1339 0.1827 1.326 0.2013 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3413 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.0427 1.616 0.4693 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.8139 0.5307 ;
        RECT 0.8139 0.4933 0.91 0.5307 ;
        RECT 0.91 0.4933 0.974 0.5307 ;
        RECT 0.974 0.4933 1.102 0.5307 ;
        RECT 1.102 0.4933 1.188 0.5307 ;
        RECT 1.188 0.4933 1.488 0.5307 ;
        RECT 1.488 0.4933 1.674 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.674 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.14 1.1339 0.1587 ;
        RECT 0.082 0.3533 1.1339 0.372 ;
      LAYER MINT1 ;
        RECT 0.146 0.14 1.1339 0.1587 ;
        RECT 0.082 0.3533 1.1339 0.372 ;
      LAYER M1 ;
        RECT 0.178 0.048 0.206 0.4639 ;
        RECT 0.306 0.048 0.334 0.4639 ;
        RECT 0.53 0.4153 0.8139 0.454 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.292 ;
        RECT 0.434 0.292 0.462 0.4467 ;
        RECT 0.462 0.0679 0.8 0.0867 ;
        RECT 0.8 0.0679 0.828 0.0867 ;
        RECT 0.8 0.0867 0.828 0.292 ;
        RECT 0.576 0.22 0.604 0.3373 ;
        RECT 0.576 0.3373 0.604 0.356 ;
        RECT 0.604 0.3373 0.882 0.356 ;
        RECT 0.882 0.048 0.91 0.22 ;
        RECT 0.882 0.22 0.91 0.3373 ;
        RECT 0.882 0.3373 0.91 0.356 ;
        RECT 0.882 0.356 0.91 0.448 ;
        RECT 1.01 0.0679 1.038 0.0867 ;
        RECT 1.01 0.0867 1.038 0.244 ;
        RECT 1.01 0.244 1.038 0.4467 ;
        RECT 1.038 0.0679 1.335 0.0867 ;
        RECT 1.335 0.0679 1.363 0.0867 ;
        RECT 1.335 0.0867 1.363 0.244 ;
        RECT 1.224 0.2627 1.252 0.4253 ;
        RECT 1.224 0.4253 1.252 0.444 ;
        RECT 1.252 0.4253 1.458 0.444 ;
        RECT 1.458 0.048 1.486 0.088 ;
        RECT 1.458 0.088 1.486 0.2627 ;
        RECT 1.458 0.2627 1.486 0.4253 ;
        RECT 1.458 0.4253 1.486 0.444 ;
        RECT 1.486 0.088 1.488 0.2627 ;
        RECT 1.486 0.2627 1.488 0.4253 ;
        RECT 1.486 0.4253 1.488 0.444 ;
        RECT 0.048 0.0567 0.08 0.0939 ;
        RECT 0.048 0.0939 0.08 0.1127 ;
        RECT 0.048 0.3779 0.08 0.404 ;
        RECT 0.048 0.404 0.08 0.4573 ;
        RECT 0.08 0.0939 0.114 0.1127 ;
        RECT 0.08 0.3779 0.114 0.404 ;
        RECT 0.114 0.0939 0.1419 0.1127 ;
        RECT 0.114 0.1127 0.1419 0.3779 ;
        RECT 0.114 0.3779 0.1419 0.404 ;
        RECT 0.37 0.1293 0.398 0.3293 ;
        RECT 0.498 0.268 0.526 0.3827 ;
        RECT 0.526 0.1293 0.558 0.196 ;
        RECT 0.736 0.172 0.764 0.292 ;
        RECT 0.946 0.1827 0.974 0.3853 ;
        RECT 1.074 0.1159 1.102 0.2113 ;
        RECT 1.074 0.3067 1.102 0.4147 ;
        RECT 1.156 0.1107 1.188 0.4573 ;
        RECT 1.266 0.1159 1.294 0.212 ;
      LAYER V1 ;
        RECT 0.114 0.3533 0.1419 0.372 ;
        RECT 0.178 0.14 0.206 0.1587 ;
        RECT 0.37 0.14 0.398 0.1587 ;
        RECT 0.498 0.3533 0.526 0.372 ;
        RECT 0.53 0.14 0.558 0.1587 ;
        RECT 0.736 0.1827 0.764 0.2013 ;
        RECT 0.946 0.3533 0.974 0.372 ;
        RECT 1.074 0.14 1.102 0.1587 ;
        RECT 1.074 0.3533 1.102 0.372 ;
        RECT 1.266 0.1827 1.294 0.2013 ;
      LAYER M1 ;
        RECT 0.178 0.048 0.206 0.4639 ;
        RECT 0.306 0.048 0.334 0.4639 ;
        RECT 0.53 0.4153 0.8139 0.454 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.292 ;
        RECT 0.434 0.292 0.462 0.4467 ;
        RECT 0.462 0.0679 0.8 0.0867 ;
        RECT 0.8 0.0679 0.828 0.0867 ;
        RECT 0.8 0.0867 0.828 0.292 ;
        RECT 0.576 0.22 0.604 0.3373 ;
        RECT 0.576 0.3373 0.604 0.356 ;
        RECT 0.604 0.3373 0.882 0.356 ;
        RECT 0.882 0.048 0.91 0.22 ;
        RECT 0.882 0.22 0.91 0.3373 ;
        RECT 0.882 0.3373 0.91 0.356 ;
        RECT 0.882 0.356 0.91 0.448 ;
        RECT 1.01 0.0679 1.038 0.0867 ;
        RECT 1.01 0.0867 1.038 0.244 ;
        RECT 1.01 0.244 1.038 0.4467 ;
        RECT 1.038 0.0679 1.335 0.0867 ;
        RECT 1.335 0.0679 1.363 0.0867 ;
        RECT 1.335 0.0867 1.363 0.244 ;
        RECT 1.224 0.2627 1.252 0.4253 ;
        RECT 1.224 0.4253 1.252 0.444 ;
        RECT 1.252 0.4253 1.458 0.444 ;
        RECT 1.458 0.048 1.486 0.088 ;
        RECT 1.458 0.088 1.486 0.2627 ;
        RECT 1.458 0.2627 1.486 0.4253 ;
        RECT 1.458 0.4253 1.486 0.444 ;
        RECT 1.486 0.088 1.488 0.2627 ;
        RECT 1.486 0.2627 1.488 0.4253 ;
        RECT 1.486 0.4253 1.488 0.444 ;
        RECT 0.048 0.0567 0.08 0.0939 ;
        RECT 0.048 0.0939 0.08 0.1127 ;
        RECT 0.048 0.3779 0.08 0.404 ;
        RECT 0.048 0.404 0.08 0.4573 ;
        RECT 0.08 0.0939 0.114 0.1127 ;
        RECT 0.08 0.3779 0.114 0.404 ;
        RECT 0.114 0.0939 0.1419 0.1127 ;
        RECT 0.114 0.1127 0.1419 0.3779 ;
        RECT 0.114 0.3779 0.1419 0.404 ;
        RECT 0.37 0.1293 0.398 0.3293 ;
        RECT 0.498 0.268 0.526 0.3827 ;
        RECT 0.526 0.1293 0.558 0.196 ;
        RECT 0.736 0.172 0.764 0.292 ;
        RECT 0.946 0.1827 0.974 0.3853 ;
        RECT 1.074 0.1159 1.102 0.2113 ;
        RECT 1.074 0.3067 1.102 0.4147 ;
        RECT 1.156 0.1107 1.188 0.4573 ;
        RECT 1.266 0.1159 1.294 0.212 ;
  END
END DFFRNQ_X1_8T

MACRO DFFSNQ_X1_8T
  CLASS core ;
  FOREIGN DFFSNQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.3507 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.722 0.1827 1.1339 0.2013 ;
        RECT 1.1339 0.1827 1.326 0.2013 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3413 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.0427 1.616 0.4693 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.554 0.5307 ;
        RECT 0.554 0.4933 0.91 0.5307 ;
        RECT 0.91 0.4933 0.974 0.5307 ;
        RECT 0.974 0.4933 1.106 0.5307 ;
        RECT 1.106 0.4933 1.3899 0.5307 ;
        RECT 1.3899 0.4933 1.488 0.5307 ;
        RECT 1.488 0.4933 1.674 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.674 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.14 1.1339 0.1587 ;
        RECT 0.082 0.3533 1.1339 0.372 ;
      LAYER MINT1 ;
        RECT 0.146 0.14 1.1339 0.1587 ;
        RECT 0.082 0.3533 1.1339 0.372 ;
      LAYER M1 ;
        RECT 0.178 0.048 0.206 0.4639 ;
        RECT 0.306 0.048 0.334 0.4639 ;
        RECT 0.434 0.0813 0.462 0.1 ;
        RECT 0.434 0.1 0.462 0.244 ;
        RECT 0.434 0.244 0.462 0.4467 ;
        RECT 0.462 0.0813 0.8179 0.1 ;
        RECT 0.8179 0.0813 0.846 0.1 ;
        RECT 0.8179 0.1 0.846 0.244 ;
        RECT 0.946 0.1827 0.974 0.3827 ;
        RECT 1.074 0.1293 1.106 0.2167 ;
        RECT 1.074 0.262 1.106 0.396 ;
        RECT 1.266 0.124 1.294 0.212 ;
        RECT 1.202 0.2627 1.23 0.3827 ;
        RECT 1.202 0.3827 1.23 0.4013 ;
        RECT 1.23 0.3827 1.458 0.4013 ;
        RECT 1.458 0.048 1.486 0.088 ;
        RECT 1.458 0.088 1.486 0.2627 ;
        RECT 1.458 0.2627 1.486 0.3827 ;
        RECT 1.458 0.3827 1.486 0.4013 ;
        RECT 1.486 0.088 1.488 0.2627 ;
        RECT 1.486 0.2627 1.488 0.3827 ;
        RECT 1.486 0.3827 1.488 0.4013 ;
        RECT 0.045 0.0547 0.048 0.092 ;
        RECT 0.045 0.092 0.048 0.118 ;
        RECT 0.048 0.0547 0.08 0.092 ;
        RECT 0.048 0.092 0.08 0.118 ;
        RECT 0.048 0.3779 0.08 0.404 ;
        RECT 0.048 0.404 0.08 0.4573 ;
        RECT 0.08 0.0547 0.083 0.092 ;
        RECT 0.08 0.092 0.083 0.118 ;
        RECT 0.08 0.3779 0.083 0.404 ;
        RECT 0.083 0.092 0.114 0.118 ;
        RECT 0.083 0.3779 0.114 0.404 ;
        RECT 0.114 0.092 0.1419 0.118 ;
        RECT 0.114 0.118 0.1419 0.3779 ;
        RECT 0.114 0.3779 0.1419 0.404 ;
        RECT 0.37 0.1293 0.398 0.3293 ;
        RECT 0.498 0.268 0.526 0.3933 ;
        RECT 0.526 0.1293 0.554 0.2033 ;
        RECT 0.754 0.172 0.782 0.244 ;
        RECT 0.608 0.1827 0.636 0.3827 ;
        RECT 0.608 0.3827 0.636 0.4013 ;
        RECT 0.636 0.3827 0.878 0.4013 ;
        RECT 0.878 0.3827 0.882 0.4013 ;
        RECT 0.878 0.4013 0.882 0.4573 ;
        RECT 0.882 0.064 0.91 0.1827 ;
        RECT 0.882 0.1827 0.91 0.3827 ;
        RECT 0.882 0.3827 0.91 0.4013 ;
        RECT 0.882 0.4013 0.91 0.4573 ;
        RECT 1.01 0.076 1.038 0.0946 ;
        RECT 1.01 0.0946 1.038 0.244 ;
        RECT 1.01 0.244 1.038 0.448 ;
        RECT 1.038 0.076 1.352 0.0946 ;
        RECT 1.352 0.076 1.3799 0.0946 ;
        RECT 1.352 0.0946 1.3799 0.244 ;
        RECT 1.106 0.4253 1.3899 0.444 ;
      LAYER V1 ;
        RECT 0.114 0.3533 0.1419 0.372 ;
        RECT 0.178 0.14 0.206 0.1587 ;
        RECT 0.37 0.14 0.398 0.1587 ;
        RECT 0.498 0.3533 0.526 0.372 ;
        RECT 0.526 0.14 0.554 0.1587 ;
        RECT 0.754 0.1827 0.782 0.2013 ;
        RECT 0.946 0.3533 0.974 0.372 ;
        RECT 1.074 0.14 1.102 0.1587 ;
        RECT 1.074 0.3533 1.102 0.372 ;
        RECT 1.266 0.1827 1.294 0.2013 ;
      LAYER M1 ;
        RECT 0.178 0.048 0.206 0.4639 ;
        RECT 0.306 0.048 0.334 0.4639 ;
        RECT 0.434 0.0813 0.462 0.1 ;
        RECT 0.434 0.1 0.462 0.244 ;
        RECT 0.434 0.244 0.462 0.4467 ;
        RECT 0.462 0.0813 0.8179 0.1 ;
        RECT 0.8179 0.0813 0.846 0.1 ;
        RECT 0.8179 0.1 0.846 0.244 ;
        RECT 0.946 0.1827 0.974 0.3827 ;
        RECT 1.074 0.1293 1.106 0.2167 ;
        RECT 1.074 0.262 1.106 0.396 ;
        RECT 1.266 0.124 1.294 0.212 ;
        RECT 1.202 0.2627 1.23 0.3827 ;
        RECT 1.202 0.3827 1.23 0.4013 ;
        RECT 1.23 0.3827 1.458 0.4013 ;
        RECT 1.458 0.048 1.486 0.088 ;
        RECT 1.458 0.088 1.486 0.2627 ;
        RECT 1.458 0.2627 1.486 0.3827 ;
        RECT 1.458 0.3827 1.486 0.4013 ;
        RECT 1.486 0.088 1.488 0.2627 ;
        RECT 1.486 0.2627 1.488 0.3827 ;
        RECT 1.486 0.3827 1.488 0.4013 ;
        RECT 0.045 0.0547 0.048 0.092 ;
        RECT 0.045 0.092 0.048 0.118 ;
        RECT 0.048 0.0547 0.08 0.092 ;
        RECT 0.048 0.092 0.08 0.118 ;
        RECT 0.048 0.3779 0.08 0.404 ;
        RECT 0.048 0.404 0.08 0.4573 ;
        RECT 0.08 0.0547 0.083 0.092 ;
        RECT 0.08 0.092 0.083 0.118 ;
        RECT 0.08 0.3779 0.083 0.404 ;
        RECT 0.083 0.092 0.114 0.118 ;
        RECT 0.083 0.3779 0.114 0.404 ;
        RECT 0.114 0.092 0.1419 0.118 ;
        RECT 0.114 0.118 0.1419 0.3779 ;
        RECT 0.114 0.3779 0.1419 0.404 ;
        RECT 0.37 0.1293 0.398 0.3293 ;
        RECT 0.498 0.268 0.526 0.3933 ;
        RECT 0.526 0.1293 0.554 0.2033 ;
        RECT 0.754 0.172 0.782 0.244 ;
        RECT 0.608 0.1827 0.636 0.3827 ;
        RECT 0.608 0.3827 0.636 0.4013 ;
        RECT 0.636 0.3827 0.878 0.4013 ;
        RECT 0.878 0.3827 0.882 0.4013 ;
        RECT 0.878 0.4013 0.882 0.4573 ;
        RECT 0.882 0.064 0.91 0.1827 ;
        RECT 0.882 0.1827 0.91 0.3827 ;
        RECT 0.882 0.3827 0.91 0.4013 ;
        RECT 0.882 0.4013 0.91 0.4573 ;
        RECT 1.01 0.076 1.038 0.0946 ;
        RECT 1.01 0.0946 1.038 0.244 ;
        RECT 1.01 0.244 1.038 0.448 ;
        RECT 1.038 0.076 1.352 0.0946 ;
        RECT 1.352 0.076 1.3799 0.0946 ;
        RECT 1.352 0.0946 1.3799 0.244 ;
        RECT 1.106 0.4253 1.3899 0.444 ;
  END
END DFFSNQ_X1_8T

MACRO FA_X1_8T
  CLASS core ;
  FOREIGN FA_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.536 BY 0.512 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.21 0.3107 1.098 0.3293 ;
      LAYER V1 ;
        RECT 0.656 0.3107 0.684 0.3293 ;
        RECT 1.038 0.3107 1.066 0.3293 ;
      LAYER M1 ;
        RECT 0.656 0.268 0.684 0.3507 ;
        RECT 1.038 0.1827 1.074 0.3507 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.1827 0.1827 0.789 0.2013 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.146 0.14 1.262 0.1587 ;
      LAYER V1 ;
        RECT 0.178 0.14 0.206 0.1587 ;
        RECT 0.58 0.14 0.608 0.1587 ;
        RECT 1.202 0.14 1.23 0.1587 ;
      LAYER M1 ;
        RECT 0.178 0.1293 0.206 0.3933 ;
        RECT 0.58 0.1293 0.608 0.244 ;
        RECT 1.202 0.1187 1.23 0.244 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.458 0.076 1.486 0.436 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8179 0.138 0.846 0.4267 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.656 0.5307 ;
        RECT 0.656 0.4933 0.767 0.5307 ;
        RECT 0.767 0.4933 1.038 0.5307 ;
        RECT 1.038 0.4933 1.084 0.5307 ;
        RECT 1.084 0.4933 1.166 0.5307 ;
        RECT 1.166 0.4933 1.289 0.5307 ;
        RECT 1.289 0.4933 1.358 0.5307 ;
        RECT 1.358 0.4933 1.546 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.546 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.082 0.268 1.321 0.2867 ;
        RECT 0.402 0.2253 1.3899 0.244 ;
      LAYER MINT1 ;
        RECT 0.082 0.268 1.321 0.2867 ;
        RECT 0.402 0.2253 1.3899 0.244 ;
      LAYER M1 ;
        RECT 0.027 0.1187 0.065 0.2253 ;
        RECT 0.027 0.2253 0.065 0.244 ;
        RECT 0.065 0.2253 0.103 0.244 ;
        RECT 0.103 0.2253 0.1419 0.244 ;
        RECT 0.103 0.244 0.1419 0.308 ;
        RECT 0.242 0.1827 0.27 0.3933 ;
        RECT 0.424 0.1827 0.462 0.338 ;
        RECT 0.37 0.0647 0.618 0.09 ;
        RECT 0.37 0.3833 0.402 0.402 ;
        RECT 0.37 0.402 0.402 0.4653 ;
        RECT 0.402 0.3833 0.624 0.402 ;
        RECT 0.624 0.3833 0.656 0.402 ;
        RECT 0.624 0.402 0.656 0.4653 ;
        RECT 0.624 0.4653 0.656 0.4693 ;
        RECT 0.729 0.1627 0.767 0.3093 ;
        RECT 0.882 0.1293 0.91 0.244 ;
        RECT 0.882 0.3747 0.91 0.3933 ;
        RECT 0.882 0.3933 0.91 0.4639 ;
        RECT 0.91 0.3747 1.01 0.3933 ;
        RECT 1.01 0.3747 1.038 0.3933 ;
        RECT 1.01 0.3933 1.038 0.4639 ;
        RECT 1.1379 0.048 1.166 0.4639 ;
        RECT 1.2609 0.2573 1.289 0.3933 ;
        RECT 0.306 0.064 0.334 0.448 ;
        RECT 0.498 0.1827 0.526 0.338 ;
        RECT 0.946 0.1827 0.984 0.3293 ;
        RECT 0.846 0.0667 1.084 0.066732 ;
        RECT 1.33 0.1827 1.358 0.3507 ;
      LAYER V1 ;
        RECT 0.114 0.268 0.1419 0.2867 ;
        RECT 0.242 0.3107 0.27 0.3293 ;
        RECT 0.306 0.1827 0.334 0.2013 ;
        RECT 0.434 0.2253 0.462 0.244 ;
        RECT 0.498 0.268 0.526 0.2867 ;
        RECT 0.729 0.1827 0.757 0.2013 ;
        RECT 0.882 0.14 0.91 0.1587 ;
        RECT 0.956 0.268 0.984 0.2867 ;
        RECT 1.1379 0.2253 1.166 0.244 ;
        RECT 1.2609 0.268 1.289 0.2867 ;
        RECT 1.33 0.2253 1.358 0.244 ;
      LAYER M1 ;
        RECT 0.027 0.1187 0.065 0.2253 ;
        RECT 0.027 0.2253 0.065 0.244 ;
        RECT 0.065 0.2253 0.103 0.244 ;
        RECT 0.103 0.2253 0.1419 0.244 ;
        RECT 0.103 0.244 0.1419 0.308 ;
        RECT 0.242 0.1827 0.27 0.3933 ;
        RECT 0.424 0.1827 0.462 0.338 ;
        RECT 0.37 0.0647 0.618 0.09 ;
        RECT 0.37 0.3833 0.402 0.402 ;
        RECT 0.37 0.402 0.402 0.4653 ;
        RECT 0.402 0.3833 0.624 0.402 ;
        RECT 0.624 0.3833 0.656 0.402 ;
        RECT 0.624 0.402 0.656 0.4653 ;
        RECT 0.624 0.4653 0.656 0.4693 ;
        RECT 0.729 0.1627 0.767 0.3093 ;
        RECT 0.882 0.1293 0.91 0.244 ;
        RECT 0.882 0.3747 0.91 0.3933 ;
        RECT 0.882 0.3933 0.91 0.4639 ;
        RECT 0.91 0.3747 1.01 0.3933 ;
        RECT 1.01 0.3747 1.038 0.3933 ;
        RECT 1.01 0.3933 1.038 0.4639 ;
        RECT 1.1379 0.048 1.166 0.4639 ;
        RECT 1.2609 0.2573 1.289 0.3933 ;
        RECT 0.306 0.064 0.334 0.448 ;
        RECT 0.498 0.1827 0.526 0.338 ;
        RECT 0.946 0.1827 0.984 0.3293 ;
        RECT 0.846 0.0667 1.084 0.066732 ;
        RECT 1.33 0.1827 1.358 0.3507 ;
  END
END FA_X1_8T

MACRO FILLTIE_8T
  CLASS core ;
  FOREIGN FILLTIE_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.578 BY 0.512 ;
  OBS
      LAYER M1 ;
        RECT -0.01 -0.0187 0.588 0.0187 ;
        RECT -0.01 0.4933 0.588 0.5307 ;
      LAYER M1 ;
        RECT -0.01 -0.0187 0.588 0.0187 ;
        RECT -0.01 0.4933 0.588 0.5307 ;
  END
END FILLTIE_8T

MACRO FILL_X1_8T
  CLASS core ;
  FOREIGN FILL_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.128 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.138 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.138 0.0187 ;
    END
  END VSS
END FILL_X1_8T

MACRO FILL_X2_8T
  CLASS core ;
  FOREIGN FILL_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.202 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.202 0.0187 ;
    END
  END VSS
END FILL_X2_8T

MACRO FILL_X4_8T
  CLASS core ;
  FOREIGN FILL_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
END FILL_X4_8T

MACRO FILL_X8_8T
  CLASS core ;
  FOREIGN FILL_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
END FILL_X8_8T

MACRO FILL_X16_8T
  CLASS core ;
  FOREIGN FILL_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.088 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.098 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.098 0.0187 ;
    END
  END VSS
END FILL_X16_8T

MACRO HA_X1_8T
  CLASS core ;
  FOREIGN HA_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.832 BY 0.512 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1827 0.27 0.3707 ;
        RECT 0.242 0.3707 0.27 0.3893 ;
        RECT 0.27 0.3707 0.434 0.3893 ;
        RECT 0.434 0.1827 0.462 0.3707 ;
        RECT 0.434 0.3707 0.462 0.3893 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.1707 0.334 0.3413 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0547 0.078 0.4253 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.754 0.12 0.782 0.4253 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.596 0.5307 ;
        RECT 0.596 0.4933 0.66 0.5307 ;
        RECT 0.66 0.4933 0.842 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.842 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.338 0.0679 0.622 0.0867 ;
        RECT 0.406 0.1227 0.498 0.144 ;
        RECT 0.498 0.1227 0.53 0.144 ;
        RECT 0.498 0.144 0.53 0.308 ;
        RECT 0.498 0.308 0.53 0.4013 ;
        RECT 0.53 0.1227 0.632 0.144 ;
        RECT 0.632 0.1227 0.66 0.144 ;
        RECT 0.632 0.144 0.66 0.308 ;
        RECT 0.114 0.1107 0.1419 0.132 ;
        RECT 0.114 0.132 0.1419 0.1827 ;
        RECT 0.114 0.1827 0.1419 0.4253 ;
        RECT 0.114 0.4253 0.1419 0.444 ;
        RECT 0.1419 0.1107 0.37 0.132 ;
        RECT 0.1419 0.4253 0.37 0.444 ;
        RECT 0.37 0.4253 0.5659 0.444 ;
        RECT 0.5659 0.1827 0.596 0.4253 ;
        RECT 0.5659 0.4253 0.596 0.444 ;
      LAYER M1 ;
        RECT 0.338 0.0679 0.622 0.0867 ;
        RECT 0.406 0.1227 0.498 0.144 ;
        RECT 0.498 0.1227 0.53 0.144 ;
        RECT 0.498 0.144 0.53 0.308 ;
        RECT 0.498 0.308 0.53 0.4013 ;
        RECT 0.53 0.1227 0.632 0.144 ;
        RECT 0.632 0.1227 0.66 0.144 ;
        RECT 0.632 0.144 0.66 0.308 ;
        RECT 0.114 0.1107 0.1419 0.132 ;
        RECT 0.114 0.132 0.1419 0.1827 ;
        RECT 0.114 0.1827 0.1419 0.4253 ;
        RECT 0.114 0.4253 0.1419 0.444 ;
        RECT 0.1419 0.1107 0.37 0.132 ;
        RECT 0.1419 0.4253 0.37 0.444 ;
        RECT 0.37 0.4253 0.5659 0.444 ;
        RECT 0.5659 0.1827 0.596 0.4253 ;
        RECT 0.5659 0.4253 0.596 0.444 ;
  END
END HA_X1_8T

MACRO INV_X1_8T
  CLASS core ;
  FOREIGN INV_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.076 0.076 0.1419 0.4267 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.202 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.202 0.0187 ;
    END
  END VSS
END INV_X1_8T

MACRO INV_X2_8T
  CLASS core ;
  FOREIGN INV_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0867 0.1419 0.384 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.266 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.266 0.0187 ;
    END
  END VSS
END INV_X2_8T

MACRO INV_X4_8T
  CLASS core ;
  FOREIGN INV_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.1707 0.08 0.2453 ;
        RECT 0.048 0.2453 0.08 0.264 ;
        RECT 0.048 0.264 0.08 0.3413 ;
        RECT 0.08 0.2453 0.238 0.264 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.0946 0.059 0.1333 ;
        RECT 0.059 0.0946 0.306 0.1333 ;
        RECT 0.059 0.3786 0.306 0.4173 ;
        RECT 0.306 0.0946 0.334 0.1333 ;
        RECT 0.306 0.1333 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4173 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END INV_X4_8T

MACRO INV_X8_8T
  CLASS core ;
  FOREIGN INV_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1293 0.1419 0.264 ;
        RECT 0.114 0.264 0.1419 0.3033 ;
        RECT 0.114 0.3033 0.1419 0.384 ;
        RECT 0.1419 0.264 0.462 0.3033 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.4207 0.054 0.4393 ;
        RECT 0.054 0.0733 0.557 0.092 ;
        RECT 0.054 0.4207 0.557 0.4393 ;
        RECT 0.557 0.0733 0.595 0.092 ;
        RECT 0.557 0.092 0.595 0.4207 ;
        RECT 0.557 0.4207 0.595 0.4393 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.65 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.65 0.0187 ;
    END
  END VSS
END INV_X8_8T

MACRO INV_X12_8T
  CLASS core ;
  FOREIGN INV_X12_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.128 0.1419 0.2453 ;
        RECT 0.114 0.2453 0.1419 0.264 ;
        RECT 0.114 0.264 0.1419 0.384 ;
        RECT 0.1419 0.2453 0.686 0.264 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.0679 0.8129 0.0867 ;
        RECT 0.054 0.424 0.8129 0.4453 ;
        RECT 0.8129 0.0679 0.851 0.0867 ;
        RECT 0.8129 0.0867 0.851 0.424 ;
        RECT 0.8129 0.424 0.851 0.4453 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.906 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.906 0.0187 ;
    END
  END VSS
END INV_X12_8T

MACRO INV_X16_8T
  CLASS core ;
  FOREIGN INV_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.152 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.2467 ;
        RECT 0.05 0.2467 0.078 0.2653 ;
        RECT 0.05 0.2653 0.078 0.3753 ;
        RECT 0.078 0.2467 0.942 0.2653 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.07 0.5307 ;
        RECT 1.07 0.4933 1.162 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.162 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.0667 1.038 0.066732 ;
        RECT 0.054 0.4147 1.038 0.454 ;
        RECT 1.038 0.0667 1.07 0.066732 ;
        RECT 1.038 0.088 1.07 0.4147 ;
        RECT 1.038 0.4147 1.07 0.454 ;
      LAYER M1 ;
        RECT 0.054 0.0667 1.038 0.066732 ;
        RECT 0.054 0.4147 1.038 0.454 ;
        RECT 1.038 0.0667 1.07 0.066732 ;
        RECT 1.038 0.088 1.07 0.4147 ;
        RECT 1.038 0.4147 1.07 0.454 ;
  END
END INV_X16_8T

MACRO LHQ_X1_8T
  CLASS core ;
  FOREIGN LHQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1067 0.27 0.3413 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3413 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8179 0.0867 0.846 0.4253 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.782 0.5307 ;
        RECT 0.782 0.4933 0.906 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.906 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.3707 0.05 0.3893 ;
        RECT 0.048 0.3893 0.05 0.4693 ;
        RECT 0.05 0.0427 0.078 0.0613 ;
        RECT 0.05 0.0613 0.078 0.1227 ;
        RECT 0.05 0.1227 0.078 0.1413 ;
        RECT 0.05 0.3707 0.078 0.3893 ;
        RECT 0.05 0.3893 0.078 0.4693 ;
        RECT 0.078 0.0427 0.08 0.0613 ;
        RECT 0.078 0.1227 0.08 0.1413 ;
        RECT 0.078 0.3707 0.08 0.3893 ;
        RECT 0.078 0.3893 0.08 0.4693 ;
        RECT 0.08 0.0427 0.114 0.0613 ;
        RECT 0.08 0.1227 0.114 0.1413 ;
        RECT 0.08 0.3707 0.114 0.3893 ;
        RECT 0.114 0.0427 0.1419 0.0613 ;
        RECT 0.114 0.1227 0.1419 0.1413 ;
        RECT 0.114 0.1413 0.1419 0.2147 ;
        RECT 0.114 0.2147 0.1419 0.2333 ;
        RECT 0.114 0.2333 0.1419 0.276 ;
        RECT 0.114 0.276 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.0427 0.324 0.0613 ;
        RECT 0.324 0.0427 0.352 0.0613 ;
        RECT 0.324 0.0613 0.352 0.1227 ;
        RECT 0.324 0.1227 0.352 0.1413 ;
        RECT 0.324 0.1413 0.352 0.2147 ;
        RECT 0.324 0.2147 0.23332 0.2333 ;
        RECT 0.23332 0.2147 0.37 0.2333 ;
        RECT 0.37 0.2147 0.398 0.2333 ;
        RECT 0.37 0.2333 0.398 0.276 ;
        RECT 0.53 0.076 0.558 0.0946 ;
        RECT 0.53 0.0946 0.558 0.3293 ;
        RECT 0.558 0.076 0.6899 0.0946 ;
        RECT 0.6899 0.076 0.718 0.0946 ;
        RECT 0.6899 0.0946 0.718 0.3293 ;
        RECT 0.6899 0.3293 0.718 0.3953 ;
        RECT 0.178 0.0907 0.206 0.3067 ;
        RECT 0.178 0.3067 0.206 0.3707 ;
        RECT 0.178 0.3707 0.206 0.3893 ;
        RECT 0.206 0.3707 0.306 0.3893 ;
        RECT 0.306 0.3067 0.34 0.3707 ;
        RECT 0.306 0.3707 0.34 0.3893 ;
        RECT 0.274 0.4253 0.388 0.444 ;
        RECT 0.388 0.076 0.466 0.1153 ;
        RECT 0.388 0.4253 0.466 0.444 ;
        RECT 0.466 0.076 0.494 0.1153 ;
        RECT 0.466 0.1153 0.494 0.204 ;
        RECT 0.466 0.204 0.494 0.4247 ;
        RECT 0.466 0.4247 0.494 0.4253 ;
        RECT 0.466 0.4253 0.494 0.444 ;
        RECT 0.494 0.4247 0.754 0.4253 ;
        RECT 0.494 0.4253 0.754 0.444 ;
        RECT 0.754 0.204 0.782 0.4247 ;
        RECT 0.754 0.4247 0.782 0.4253 ;
        RECT 0.754 0.4253 0.782 0.444 ;
      LAYER M1 ;
        RECT 0.048 0.3707 0.05 0.3893 ;
        RECT 0.048 0.3893 0.05 0.4693 ;
        RECT 0.05 0.0427 0.078 0.0613 ;
        RECT 0.05 0.0613 0.078 0.1227 ;
        RECT 0.05 0.1227 0.078 0.1413 ;
        RECT 0.05 0.3707 0.078 0.3893 ;
        RECT 0.05 0.3893 0.078 0.4693 ;
        RECT 0.078 0.0427 0.08 0.0613 ;
        RECT 0.078 0.1227 0.08 0.1413 ;
        RECT 0.078 0.3707 0.08 0.3893 ;
        RECT 0.078 0.3893 0.08 0.4693 ;
        RECT 0.08 0.0427 0.114 0.0613 ;
        RECT 0.08 0.1227 0.114 0.1413 ;
        RECT 0.08 0.3707 0.114 0.3893 ;
        RECT 0.114 0.0427 0.1419 0.0613 ;
        RECT 0.114 0.1227 0.1419 0.1413 ;
        RECT 0.114 0.1413 0.1419 0.2147 ;
        RECT 0.114 0.2147 0.1419 0.2333 ;
        RECT 0.114 0.2333 0.1419 0.276 ;
        RECT 0.114 0.276 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.0427 0.324 0.0613 ;
        RECT 0.324 0.0427 0.352 0.0613 ;
        RECT 0.324 0.0613 0.352 0.1227 ;
        RECT 0.324 0.1227 0.352 0.1413 ;
        RECT 0.324 0.1413 0.352 0.2147 ;
        RECT 0.324 0.2147 0.23332 0.2333 ;
        RECT 0.23332 0.2147 0.37 0.2333 ;
        RECT 0.37 0.2147 0.398 0.2333 ;
        RECT 0.37 0.2333 0.398 0.276 ;
        RECT 0.53 0.076 0.558 0.0946 ;
        RECT 0.53 0.0946 0.558 0.3293 ;
        RECT 0.558 0.076 0.6899 0.0946 ;
        RECT 0.6899 0.076 0.718 0.0946 ;
        RECT 0.6899 0.0946 0.718 0.3293 ;
        RECT 0.6899 0.3293 0.718 0.3953 ;
        RECT 0.178 0.0907 0.206 0.3067 ;
        RECT 0.178 0.3067 0.206 0.3707 ;
        RECT 0.178 0.3707 0.206 0.3893 ;
        RECT 0.206 0.3707 0.306 0.3893 ;
        RECT 0.306 0.3067 0.34 0.3707 ;
        RECT 0.306 0.3707 0.34 0.3893 ;
        RECT 0.274 0.4253 0.388 0.444 ;
        RECT 0.388 0.076 0.466 0.1153 ;
        RECT 0.388 0.4253 0.466 0.444 ;
        RECT 0.466 0.076 0.494 0.1153 ;
        RECT 0.466 0.1153 0.494 0.204 ;
        RECT 0.466 0.204 0.494 0.4247 ;
        RECT 0.466 0.4247 0.494 0.4253 ;
        RECT 0.466 0.4253 0.494 0.444 ;
        RECT 0.494 0.4247 0.754 0.4253 ;
        RECT 0.494 0.4253 0.754 0.444 ;
        RECT 0.754 0.204 0.782 0.4247 ;
        RECT 0.754 0.4247 0.782 0.4253 ;
        RECT 0.754 0.4253 0.782 0.444 ;
  END
END LHQ_X1_8T

MACRO MUX2_X1_8T
  CLASS core ;
  FOREIGN MUX2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.832 BY 0.512 ;
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.1613 0.59 0.3507 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.2987 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.118 0.4387 0.394 0.4573 ;
      LAYER V1 ;
        RECT 0.15 0.4387 0.206 0.4573 ;
      LAYER M1 ;
        RECT 0.027 0.1613 0.055 0.4387 ;
        RECT 0.027 0.4387 0.055 0.4573 ;
        RECT 0.055 0.4387 0.222 0.4573 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.6899 0.128 0.718 0.4253 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.462 0.5307 ;
        RECT 0.462 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.782 0.5307 ;
        RECT 0.782 0.4933 0.842 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.842 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.274 0.2253 0.558 0.244 ;
      LAYER MINT1 ;
        RECT 0.274 0.2253 0.558 0.244 ;
      LAYER M1 ;
        RECT 0.08 0.108 0.099 0.1267 ;
        RECT 0.099 0.108 0.157 0.1267 ;
        RECT 0.099 0.328 0.157 0.3467 ;
        RECT 0.099 0.3467 0.157 0.384 ;
        RECT 0.157 0.108 0.306 0.1267 ;
        RECT 0.157 0.328 0.306 0.3467 ;
        RECT 0.306 0.108 0.334 0.1267 ;
        RECT 0.306 0.1267 0.334 0.328 ;
        RECT 0.306 0.328 0.334 0.3467 ;
        RECT 0.29 0.4387 0.434 0.4693 ;
        RECT 0.434 0.204 0.462 0.4387 ;
        RECT 0.434 0.4387 0.462 0.4693 ;
        RECT 0.498 0.1827 0.526 0.2853 ;
        RECT 0.37 0.0579 0.398 0.0973 ;
        RECT 0.37 0.0973 0.398 0.3293 ;
        RECT 0.37 0.3293 0.398 0.4093 ;
        RECT 0.398 0.0579 0.754 0.0973 ;
        RECT 0.754 0.0579 0.782 0.0973 ;
        RECT 0.754 0.0973 0.782 0.3293 ;
      LAYER V1 ;
        RECT 0.306 0.2253 0.334 0.244 ;
        RECT 0.306 0.4387 0.362 0.4573 ;
        RECT 0.498 0.2253 0.526 0.244 ;
      LAYER M1 ;
        RECT 0.08 0.108 0.099 0.1267 ;
        RECT 0.099 0.108 0.157 0.1267 ;
        RECT 0.099 0.328 0.157 0.3467 ;
        RECT 0.099 0.3467 0.157 0.384 ;
        RECT 0.157 0.108 0.306 0.1267 ;
        RECT 0.157 0.328 0.306 0.3467 ;
        RECT 0.306 0.108 0.334 0.1267 ;
        RECT 0.306 0.1267 0.334 0.328 ;
        RECT 0.306 0.328 0.334 0.3467 ;
        RECT 0.29 0.4387 0.434 0.4693 ;
        RECT 0.434 0.204 0.462 0.4387 ;
        RECT 0.434 0.4387 0.462 0.4693 ;
        RECT 0.498 0.1827 0.526 0.2853 ;
        RECT 0.37 0.0579 0.398 0.0973 ;
        RECT 0.37 0.0973 0.398 0.3293 ;
        RECT 0.37 0.3293 0.398 0.4093 ;
        RECT 0.398 0.0579 0.754 0.0973 ;
        RECT 0.754 0.0579 0.782 0.0973 ;
        RECT 0.754 0.0973 0.782 0.3293 ;
  END
END MUX2_X1_8T

MACRO NAND2_X1_8T
  CLASS core ;
  FOREIGN NAND2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.3827 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3827 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0887 0.1419 0.128 ;
        RECT 0.114 0.128 0.1419 0.4253 ;
        RECT 0.1419 0.0887 0.176 0.128 ;
        RECT 0.176 0.0427 0.208 0.0887 ;
        RECT 0.176 0.0887 0.208 0.128 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.266 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.266 0.0187 ;
    END
  END VSS
END NAND2_X1_8T

MACRO NAND2_X2_8T
  CLASS core ;
  FOREIGN NAND2_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.15 0.206 0.3687 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1827 0.078 0.4507 ;
        RECT 0.05 0.4507 0.078 0.4693 ;
        RECT 0.078 0.4507 0.306 0.4693 ;
        RECT 0.306 0.1827 0.334 0.4507 ;
        RECT 0.306 0.4507 0.334 0.4693 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.082 0.1419 0.1207 ;
        RECT 0.114 0.1207 0.1419 0.2827 ;
        RECT 0.114 0.2827 0.1419 0.398 ;
        RECT 0.114 0.398 0.1419 0.4267 ;
        RECT 0.1419 0.082 0.242 0.1207 ;
        RECT 0.1419 0.398 0.242 0.4267 ;
        RECT 0.242 0.082 0.27 0.1207 ;
        RECT 0.242 0.2827 0.27 0.398 ;
        RECT 0.242 0.398 0.27 0.4267 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END NAND2_X2_8T

MACRO NAND3_X1_8T
  CLASS core ;
  FOREIGN NAND3_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2133 0.27 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.17 0.206 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1433 0.078 0.3827 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.07334 0.0547 0.1419 0.0733 ;
        RECT 0.07334 0.0733 0.1419 0.1707 ;
        RECT 0.114 0.1707 0.1419 0.3413 ;
        RECT 0.114 0.3413 0.1419 0.4507 ;
        RECT 0.114 0.4507 0.1419 0.4693 ;
        RECT 0.1419 0.0547 0.242 0.0733 ;
        RECT 0.1419 0.4507 0.242 0.4693 ;
        RECT 0.242 0.0427 0.304 0.0547 ;
        RECT 0.242 0.0547 0.304 0.0733 ;
        RECT 0.242 0.4507 0.304 0.4693 ;
        RECT 0.304 0.0427 0.306 0.0547 ;
        RECT 0.304 0.0547 0.306 0.0733 ;
        RECT 0.304 0.0733 0.306 0.1707 ;
        RECT 0.304 0.4507 0.306 0.4693 ;
        RECT 0.306 0.0427 0.334 0.0547 ;
        RECT 0.306 0.0547 0.334 0.0733 ;
        RECT 0.306 0.0733 0.334 0.1707 ;
        RECT 0.306 0.3413 0.334 0.4507 ;
        RECT 0.306 0.4507 0.334 0.4693 ;
        RECT 0.334 0.0427 0.336 0.0547 ;
        RECT 0.334 0.0547 0.336 0.0733 ;
        RECT 0.334 0.0733 0.336 0.1707 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END NAND3_X1_8T

MACRO NAND3_X2_8T
  CLASS core ;
  FOREIGN NAND3_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.2133 0.526 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.301 0.166 0.339 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.3413 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.027 0.3786 0.366 0.4173 ;
        RECT 0.366 0.3786 0.434 0.4173 ;
        RECT 0.434 0.124 0.462 0.3786 ;
        RECT 0.434 0.3786 0.462 0.4173 ;
        RECT 0.462 0.3786 0.494 0.4173 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.366 0.5307 ;
        RECT 0.366 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.074 0.498 0.0939 ;
        RECT 0.498 0.074 0.526 0.0939 ;
        RECT 0.498 0.0939 0.526 0.15 ;
        RECT 0.05 0.118 0.366 0.1393 ;
      LAYER M1 ;
        RECT 0.21 0.074 0.498 0.0939 ;
        RECT 0.498 0.074 0.526 0.0939 ;
        RECT 0.498 0.0939 0.526 0.15 ;
        RECT 0.05 0.118 0.366 0.1393 ;
  END
END NAND3_X2_8T

MACRO NAND4_X1_8T
  CLASS core ;
  FOREIGN NAND4_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.1707 0.398 0.3827 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1293 0.206 0.2987 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1293 0.078 0.3827 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.3413 0.1419 0.43 ;
        RECT 0.114 0.43 0.1419 0.4693 ;
        RECT 0.1419 0.43 0.306 0.4693 ;
        RECT 0.306 0.1093 0.334 0.128 ;
        RECT 0.306 0.128 0.334 0.3413 ;
        RECT 0.306 0.3413 0.334 0.43 ;
        RECT 0.306 0.43 0.334 0.4693 ;
        RECT 0.334 0.1093 0.365 0.128 ;
        RECT 0.365 0.0427 0.403 0.1093 ;
        RECT 0.365 0.1093 0.403 0.128 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
END NAND4_X1_8T

MACRO NAND4_X2_8T
  CLASS core ;
  FOREIGN NAND4_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.2387 0.594 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.2267 0.398 0.3507 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1613 0.206 0.3413 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1713 0.078 0.3413 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.37 0.144 0.384 ;
        RECT 0.112 0.384 0.144 0.4253 ;
        RECT 0.112 0.4253 0.144 0.444 ;
        RECT 0.144 0.4253 0.434 0.444 ;
        RECT 0.434 0.196 0.462 0.2147 ;
        RECT 0.434 0.2147 0.462 0.3653 ;
        RECT 0.434 0.3653 0.462 0.37 ;
        RECT 0.434 0.37 0.462 0.384 ;
        RECT 0.434 0.4253 0.462 0.444 ;
        RECT 0.462 0.196 0.562 0.2147 ;
        RECT 0.462 0.3653 0.562 0.37 ;
        RECT 0.462 0.37 0.562 0.384 ;
        RECT 0.462 0.4253 0.562 0.444 ;
        RECT 0.562 0.196 0.59 0.2147 ;
        RECT 0.562 0.3653 0.59 0.37 ;
        RECT 0.562 0.37 0.59 0.384 ;
        RECT 0.562 0.384 0.59 0.4253 ;
        RECT 0.562 0.4253 0.59 0.444 ;
        RECT 0.59 0.196 0.654 0.2147 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.656 0.5307 ;
        RECT 0.656 0.4933 0.714 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.714 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.43 0.0867 ;
        RECT 0.274 0.1533 0.624 0.172 ;
        RECT 0.624 0.0427 0.656 0.1533 ;
        RECT 0.624 0.1533 0.656 0.172 ;
        RECT 0.146 0.1107 0.494 0.1293 ;
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.43 0.0867 ;
        RECT 0.274 0.1533 0.624 0.172 ;
        RECT 0.624 0.0427 0.656 0.1533 ;
        RECT 0.624 0.1533 0.656 0.172 ;
        RECT 0.146 0.1107 0.494 0.1293 ;
  END
END NAND4_X2_8T

MACRO NOR2_X1_8T
  CLASS core ;
  FOREIGN NOR2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1293 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1293 0.078 0.3413 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0867 0.1419 0.384 ;
        RECT 0.114 0.384 0.1419 0.4233 ;
        RECT 0.1419 0.384 0.176 0.4233 ;
        RECT 0.176 0.384 0.208 0.4233 ;
        RECT 0.176 0.4233 0.208 0.4693 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.266 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.266 0.0187 ;
    END
  END VSS
END NOR2_X1_8T

MACRO NOR2_X2_8T
  CLASS core ;
  FOREIGN NOR2_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1433 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0427 0.078 0.0613 ;
        RECT 0.05 0.0613 0.078 0.3293 ;
        RECT 0.078 0.0427 0.306 0.0613 ;
        RECT 0.306 0.0427 0.334 0.0613 ;
        RECT 0.306 0.0613 0.334 0.3293 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0853 0.1419 0.104 ;
        RECT 0.114 0.104 0.1419 0.2293 ;
        RECT 0.114 0.2293 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.0853 0.176 0.104 ;
        RECT 0.1419 0.3707 0.176 0.3893 ;
        RECT 0.176 0.0853 0.208 0.104 ;
        RECT 0.176 0.3707 0.208 0.3893 ;
        RECT 0.176 0.3893 0.208 0.4267 ;
        RECT 0.208 0.0853 0.242 0.104 ;
        RECT 0.242 0.0853 0.27 0.104 ;
        RECT 0.242 0.104 0.27 0.2293 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END NOR2_X2_8T

MACRO NOR3_X1_8T
  CLASS core ;
  FOREIGN NOR3_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2133 0.27 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1293 0.206 0.3687 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1293 0.078 0.3687 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0427 0.1419 0.0613 ;
        RECT 0.114 0.0613 0.1419 0.1707 ;
        RECT 0.114 0.1707 0.1419 0.3413 ;
        RECT 0.114 0.3413 0.1419 0.4093 ;
        RECT 0.114 0.4093 0.1419 0.428 ;
        RECT 0.1419 0.0427 0.303 0.0613 ;
        RECT 0.1419 0.4093 0.303 0.428 ;
        RECT 0.303 0.0427 0.304 0.0613 ;
        RECT 0.303 0.0613 0.304 0.1707 ;
        RECT 0.303 0.4093 0.304 0.428 ;
        RECT 0.304 0.0427 0.336 0.0613 ;
        RECT 0.304 0.0613 0.336 0.1707 ;
        RECT 0.304 0.3413 0.336 0.4093 ;
        RECT 0.304 0.4093 0.336 0.428 ;
        RECT 0.304 0.428 0.336 0.4693 ;
        RECT 0.336 0.0427 0.337 0.0613 ;
        RECT 0.336 0.0613 0.337 0.1707 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END NOR3_X1_8T

MACRO NOR3_X2_8T
  CLASS core ;
  FOREIGN NOR3_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.1707 0.526 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.1707 0.334 0.342 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.346 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0859 0.1027 0.434 0.1413 ;
        RECT 0.434 0.1027 0.462 0.1413 ;
        RECT 0.434 0.1413 0.462 0.384 ;
        RECT 0.462 0.1027 0.49 0.1413 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.418 0.498 0.4367 ;
        RECT 0.498 0.344 0.526 0.418 ;
        RECT 0.498 0.418 0.526 0.4367 ;
        RECT 0.0859 0.3713 0.38 0.394 ;
      LAYER M1 ;
        RECT 0.21 0.418 0.498 0.4367 ;
        RECT 0.498 0.344 0.526 0.418 ;
        RECT 0.498 0.418 0.526 0.4367 ;
        RECT 0.0859 0.3713 0.38 0.394 ;
  END
END NOR3_X2_8T

MACRO NOR4_X1_8T
  CLASS core ;
  FOREIGN NOR4_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.1293 0.398 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1293 0.27 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.3827 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1293 0.078 0.3827 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0427 0.1419 0.0679 ;
        RECT 0.114 0.0679 0.1419 0.1433 ;
        RECT 0.1419 0.0427 0.306 0.0679 ;
        RECT 0.306 0.0427 0.334 0.0679 ;
        RECT 0.306 0.0679 0.334 0.1433 ;
        RECT 0.306 0.1433 0.334 0.384 ;
        RECT 0.306 0.384 0.334 0.4027 ;
        RECT 0.334 0.384 0.365 0.4027 ;
        RECT 0.365 0.384 0.403 0.4027 ;
        RECT 0.365 0.4027 0.403 0.4693 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
END NOR4_X1_8T

MACRO NOR4_X2_8T
  CLASS core ;
  FOREIGN NOR4_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.1707 0.594 0.2707 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.1613 0.398 0.292 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.3507 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.344 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.0679 0.144 0.0867 ;
        RECT 0.112 0.0867 0.144 0.128 ;
        RECT 0.112 0.128 0.144 0.142 ;
        RECT 0.144 0.0679 0.434 0.0867 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.128 0.462 0.142 ;
        RECT 0.434 0.142 0.462 0.1467 ;
        RECT 0.434 0.1467 0.462 0.2947 ;
        RECT 0.434 0.2947 0.462 0.3133 ;
        RECT 0.462 0.0679 0.562 0.0867 ;
        RECT 0.462 0.128 0.562 0.142 ;
        RECT 0.462 0.142 0.562 0.1467 ;
        RECT 0.462 0.2947 0.562 0.3133 ;
        RECT 0.562 0.0679 0.59 0.0867 ;
        RECT 0.562 0.0867 0.59 0.128 ;
        RECT 0.562 0.128 0.59 0.142 ;
        RECT 0.562 0.142 0.59 0.1467 ;
        RECT 0.562 0.2947 0.59 0.3133 ;
        RECT 0.59 0.2947 0.663 0.3133 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.43 0.5307 ;
        RECT 0.43 0.4933 0.494 0.5307 ;
        RECT 0.494 0.4933 0.656 0.5307 ;
        RECT 0.656 0.4933 0.714 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.714 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.3799 0.494 0.4013 ;
        RECT 0.048 0.37 0.08 0.4253 ;
        RECT 0.048 0.4253 0.08 0.444 ;
        RECT 0.08 0.4253 0.43 0.444 ;
        RECT 0.338 0.3373 0.624 0.356 ;
        RECT 0.624 0.3373 0.656 0.356 ;
        RECT 0.624 0.356 0.656 0.4573 ;
      LAYER M1 ;
        RECT 0.21 0.3799 0.494 0.4013 ;
        RECT 0.048 0.37 0.08 0.4253 ;
        RECT 0.048 0.4253 0.08 0.444 ;
        RECT 0.08 0.4253 0.43 0.444 ;
        RECT 0.338 0.3373 0.624 0.356 ;
        RECT 0.624 0.3373 0.656 0.356 ;
        RECT 0.624 0.356 0.656 0.4573 ;
  END
END NOR4_X2_8T

MACRO OAI21_X1_8T
  CLASS core ;
  FOREIGN OAI21_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.4227 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.1707 0.334 0.384 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.424 ;
        RECT 0.114 0.424 0.1419 0.4453 ;
        RECT 0.1419 0.424 0.298 0.4453 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.298 0.5307 ;
        RECT 0.298 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.0487 0.078 0.1033 ;
        RECT 0.05 0.1033 0.078 0.1247 ;
        RECT 0.078 0.1033 0.298 0.1247 ;
      LAYER M1 ;
        RECT 0.05 0.0487 0.078 0.1033 ;
        RECT 0.05 0.1033 0.078 0.1247 ;
        RECT 0.078 0.1033 0.298 0.1247 ;
  END
END OAI21_X1_8T

MACRO OAI21_X2_8T
  CLASS core ;
  FOREIGN OAI21_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.365 0.2133 0.403 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.1886 ;
        RECT 0.242 0.1886 0.27 0.3347 ;
        RECT 0.242 0.3347 0.27 0.3533 ;
        RECT 0.27 0.3347 0.498 0.3533 ;
        RECT 0.498 0.1886 0.526 0.3347 ;
        RECT 0.498 0.3347 0.526 0.3533 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.35 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.029 0.3799 0.178 0.4013 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.1853 ;
        RECT 0.178 0.1853 0.206 0.3799 ;
        RECT 0.178 0.3799 0.206 0.4013 ;
        RECT 0.206 0.1107 0.426 0.1293 ;
        RECT 0.206 0.3799 0.426 0.4013 ;
        RECT 0.426 0.1107 0.434 0.1293 ;
        RECT 0.434 0.1107 0.462 0.1293 ;
        RECT 0.434 0.1293 0.462 0.1853 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.535 0.5307 ;
        RECT 0.535 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.498 0.0867 ;
        RECT 0.498 0.0679 0.526 0.0867 ;
        RECT 0.498 0.0867 0.526 0.142 ;
        RECT 0.498 0.142 0.526 0.1433 ;
        RECT 0.146 0.4253 0.535 0.444 ;
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.498 0.0867 ;
        RECT 0.498 0.0679 0.526 0.0867 ;
        RECT 0.498 0.0867 0.526 0.142 ;
        RECT 0.498 0.142 0.526 0.1433 ;
        RECT 0.146 0.4253 0.535 0.444 ;
  END
END OAI21_X2_8T

MACRO OAI22_X1_8T
  CLASS core ;
  FOREIGN OAI22_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1327 0.27 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.186 0.398 0.384 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.128 0.206 0.3413 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.128 0.08 0.384 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1409 0.4253 0.306 0.444 ;
        RECT 0.306 0.1213 0.334 0.4253 ;
        RECT 0.306 0.4253 0.334 0.444 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.0673 0.37 0.0873 ;
        RECT 0.37 0.0673 0.398 0.0873 ;
        RECT 0.37 0.0873 0.398 0.1407 ;
      LAYER M1 ;
        RECT 0.05 0.0673 0.37 0.0873 ;
        RECT 0.37 0.0673 0.398 0.0873 ;
        RECT 0.37 0.0873 0.398 0.1407 ;
  END
END OAI22_X1_8T

MACRO OAI22_X2_8T
  CLASS core ;
  FOREIGN OAI22_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.1707 0.462 0.186 ;
        RECT 0.434 0.186 0.462 0.3107 ;
        RECT 0.434 0.3107 0.462 0.3293 ;
        RECT 0.462 0.3107 0.6899 0.3293 ;
        RECT 0.6899 0.186 0.718 0.3107 ;
        RECT 0.6899 0.3107 0.718 0.3293 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.1707 0.59 0.2653 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.1613 0.334 0.324 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1613 0.1419 0.3413 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2573 0.27 0.3533 ;
        RECT 0.242 0.3533 0.27 0.372 ;
        RECT 0.27 0.3533 0.37 0.372 ;
        RECT 0.37 0.1127 0.398 0.1313 ;
        RECT 0.37 0.1313 0.398 0.1853 ;
        RECT 0.37 0.1853 0.398 0.2573 ;
        RECT 0.37 0.2573 0.398 0.3533 ;
        RECT 0.37 0.3533 0.398 0.372 ;
        RECT 0.398 0.1127 0.626 0.1313 ;
        RECT 0.398 0.3533 0.626 0.372 ;
        RECT 0.626 0.1127 0.654 0.1313 ;
        RECT 0.626 0.1313 0.654 0.1853 ;
        RECT 0.626 0.3533 0.654 0.372 ;
        RECT 0.654 0.3533 0.6899 0.372 ;
        RECT 0.6899 0.3533 0.718 0.372 ;
        RECT 0.6899 0.372 0.718 0.448 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.362 0.5307 ;
        RECT 0.362 0.4933 0.654 0.5307 ;
        RECT 0.654 0.4933 0.718 0.5307 ;
        RECT 0.718 0.4933 0.778 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.778 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.402 0.4027 0.626 0.424 ;
        RECT 0.626 0.4027 0.654 0.424 ;
        RECT 0.626 0.424 0.654 0.4639 ;
        RECT 0.041 0.066 0.6899 0.0887 ;
        RECT 0.6899 0.066 0.718 0.0887 ;
        RECT 0.6899 0.0887 0.718 0.1407 ;
        RECT 0.05 0.408 0.362 0.4467 ;
      LAYER M1 ;
        RECT 0.402 0.4027 0.626 0.424 ;
        RECT 0.626 0.4027 0.654 0.424 ;
        RECT 0.626 0.424 0.654 0.4639 ;
        RECT 0.041 0.066 0.6899 0.0887 ;
        RECT 0.6899 0.066 0.718 0.0887 ;
        RECT 0.6899 0.0887 0.718 0.1407 ;
        RECT 0.05 0.408 0.362 0.4467 ;
  END
END OAI22_X2_8T

MACRO OR2_X1_8T
  CLASS core ;
  FOREIGN OR2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.064 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.162 0.078 0.4273 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.076 0.334 0.4267 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.0867 0.1419 0.224 ;
        RECT 0.114 0.224 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.3707 0.242 0.3893 ;
        RECT 0.242 0.224 0.27 0.3707 ;
        RECT 0.242 0.3707 0.27 0.3893 ;
      LAYER M1 ;
        RECT 0.114 0.0867 0.1419 0.224 ;
        RECT 0.114 0.224 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.3707 0.242 0.3893 ;
        RECT 0.242 0.224 0.27 0.3707 ;
        RECT 0.242 0.3707 0.27 0.3893 ;
  END
END OR2_X1_8T

MACRO OR2_X2_8T
  CLASS core ;
  FOREIGN OR2_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1613 0.1419 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3413 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.0427 0.306 0.09 ;
        RECT 0.302 0.4253 0.306 0.4693 ;
        RECT 0.306 0.0427 0.334 0.09 ;
        RECT 0.306 0.09 0.334 0.4253 ;
        RECT 0.306 0.4253 0.334 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.077 0.1027 0.146 0.1253 ;
        RECT 0.146 0.1027 0.242 0.1253 ;
        RECT 0.146 0.3867 0.242 0.4053 ;
        RECT 0.242 0.1027 0.27 0.1253 ;
        RECT 0.242 0.1253 0.27 0.3867 ;
        RECT 0.242 0.3867 0.27 0.4053 ;
      LAYER M1 ;
        RECT 0.077 0.1027 0.146 0.1253 ;
        RECT 0.146 0.1027 0.242 0.1253 ;
        RECT 0.146 0.3867 0.242 0.4053 ;
        RECT 0.242 0.1027 0.27 0.1253 ;
        RECT 0.242 0.1253 0.27 0.3867 ;
        RECT 0.242 0.3867 0.27 0.4053 ;
  END
END OR2_X2_8T

MACRO OR3_X1_8T
  CLASS core ;
  FOREIGN OR3_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.128 0.334 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.176 0.128 0.208 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.128 0.083 0.384 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.076 0.462 0.436 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.234 0.5307 ;
        RECT 0.234 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.0727 0.278 0.0913 ;
        RECT 0.278 0.0727 0.37 0.0913 ;
        RECT 0.278 0.4207 0.37 0.4487 ;
        RECT 0.37 0.0727 0.398 0.0913 ;
        RECT 0.37 0.0913 0.398 0.4207 ;
        RECT 0.37 0.4207 0.398 0.4487 ;
        RECT 0.0859 0.424 0.234 0.4453 ;
      LAYER M1 ;
        RECT 0.054 0.0727 0.278 0.0913 ;
        RECT 0.278 0.0727 0.37 0.0913 ;
        RECT 0.278 0.4207 0.37 0.4487 ;
        RECT 0.37 0.0727 0.398 0.0913 ;
        RECT 0.37 0.0913 0.398 0.4207 ;
        RECT 0.37 0.4207 0.398 0.4487 ;
        RECT 0.0859 0.424 0.234 0.4453 ;
  END
END OR3_X1_8T

MACRO OR3_X2_8T
  CLASS core ;
  FOREIGN OR3_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.17 0.1419 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3507 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.154 0.27 0.2987 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.366 0.0427 0.37 0.0867 ;
        RECT 0.366 0.424 0.37 0.4693 ;
        RECT 0.37 0.0427 0.398 0.0867 ;
        RECT 0.37 0.0867 0.398 0.424 ;
        RECT 0.37 0.424 0.398 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.302 0.5307 ;
        RECT 0.302 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.3819 0.078 0.402 ;
        RECT 0.05 0.402 0.078 0.4573 ;
        RECT 0.078 0.3819 0.302 0.402 ;
        RECT 0.06 0.1033 0.1409 0.1247 ;
        RECT 0.1409 0.1033 0.306 0.1247 ;
        RECT 0.1409 0.3367 0.306 0.358 ;
        RECT 0.306 0.1033 0.334 0.1247 ;
        RECT 0.306 0.1247 0.334 0.3367 ;
        RECT 0.306 0.3367 0.334 0.358 ;
      LAYER M1 ;
        RECT 0.05 0.3819 0.078 0.402 ;
        RECT 0.05 0.402 0.078 0.4573 ;
        RECT 0.078 0.3819 0.302 0.402 ;
        RECT 0.06 0.1033 0.1409 0.1247 ;
        RECT 0.1409 0.1033 0.306 0.1247 ;
        RECT 0.1409 0.3367 0.306 0.358 ;
        RECT 0.306 0.1033 0.334 0.1247 ;
        RECT 0.306 0.1247 0.334 0.3367 ;
        RECT 0.306 0.3367 0.334 0.358 ;
  END
END OR3_X2_8T

MACRO OR4_X1_8T
  CLASS core ;
  FOREIGN OR4_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.128 0.398 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.128 0.272 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.132 0.1419 0.384 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.076 0.526 0.4267 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.298 0.5307 ;
        RECT 0.298 0.4933 0.462 0.5307 ;
        RECT 0.462 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.0679 0.338 0.0867 ;
        RECT 0.338 0.0679 0.434 0.0867 ;
        RECT 0.338 0.42 0.434 0.4413 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.42 ;
        RECT 0.434 0.42 0.462 0.4413 ;
        RECT 0.146 0.4113 0.298 0.4367 ;
      LAYER M1 ;
        RECT 0.054 0.0679 0.338 0.0867 ;
        RECT 0.338 0.0679 0.434 0.0867 ;
        RECT 0.338 0.42 0.434 0.4413 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.42 ;
        RECT 0.434 0.42 0.462 0.4413 ;
        RECT 0.146 0.4113 0.298 0.4367 ;
  END
END OR4_X1_8T

MACRO OR4_X2_8T
  CLASS core ;
  FOREIGN OR4_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.128 0.334 0.3533 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.142 0.27 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.142 0.1419 0.384 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1273 0.078 0.384 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.496 0.0853 0.528 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.302 0.5307 ;
        RECT 0.302 0.4933 0.46 0.5307 ;
        RECT 0.46 0.4933 0.65 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.65 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.146 0.4153 0.302 0.454 ;
        RECT 0.054 0.0579 0.342 0.0967 ;
        RECT 0.342 0.0579 0.432 0.0967 ;
        RECT 0.342 0.3786 0.432 0.416 ;
        RECT 0.432 0.0579 0.46 0.0967 ;
        RECT 0.432 0.0967 0.46 0.3786 ;
        RECT 0.432 0.3786 0.46 0.416 ;
      LAYER M1 ;
        RECT 0.146 0.4153 0.302 0.454 ;
        RECT 0.054 0.0579 0.342 0.0967 ;
        RECT 0.342 0.0579 0.432 0.0967 ;
        RECT 0.342 0.3786 0.432 0.416 ;
        RECT 0.432 0.0579 0.46 0.0967 ;
        RECT 0.432 0.0967 0.46 0.3786 ;
        RECT 0.432 0.3786 0.46 0.416 ;
  END
END OR4_X2_8T

MACRO SDFFRNQ_X1_8T
  CLASS core ;
  FOREIGN SDFFRNQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.92 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.242 0.515 0.352 ;
        RECT 0.515 0.242 0.526 0.352 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.965 0.2253 1.454 0.244 ;
        RECT 1.454 0.2253 1.592 0.244 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.248 0.334 0.3813 ;
        RECT 0.306 0.3813 0.334 0.4 ;
        RECT 0.334 0.3813 0.515 0.4 ;
        RECT 0.515 0.3813 0.562 0.4 ;
        RECT 0.562 0.2093 0.59 0.248 ;
        RECT 0.562 0.248 0.59 0.3813 ;
        RECT 0.562 0.3813 0.59 0.4 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.242 0.398 0.3413 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.184 0.078 0.356 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.0427 1.872 0.4693 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.754 0.5307 ;
        RECT 0.754 0.4933 0.782 0.5307 ;
        RECT 0.782 0.4933 1.066 0.5307 ;
        RECT 1.066 0.4933 1.422 0.5307 ;
        RECT 1.422 0.4933 1.49 0.5307 ;
        RECT 1.49 0.4933 1.742 0.5307 ;
        RECT 1.742 0.4933 1.93 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.93 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.3533 1.326 0.372 ;
        RECT 0.722 0.268 1.121 0.2867 ;
        RECT 0.082 0.1827 1.454 0.2013 ;
      LAYER MINT1 ;
        RECT 0.146 0.3533 1.326 0.372 ;
        RECT 0.722 0.268 1.121 0.2867 ;
        RECT 0.082 0.1827 1.454 0.2013 ;
      LAYER M1 ;
        RECT 0.045 0.064 0.083 0.1359 ;
        RECT 0.045 0.1359 0.083 0.1547 ;
        RECT 0.045 0.4027 0.083 0.4213 ;
        RECT 0.045 0.4213 0.083 0.4586 ;
        RECT 0.083 0.1359 0.114 0.1547 ;
        RECT 0.083 0.4027 0.114 0.4213 ;
        RECT 0.114 0.1359 0.1419 0.1547 ;
        RECT 0.114 0.1547 0.1419 0.4027 ;
        RECT 0.114 0.4027 0.1419 0.4213 ;
        RECT 0.242 0.064 0.27 0.178 ;
        RECT 0.242 0.178 0.27 0.1967 ;
        RECT 0.242 0.1967 0.27 0.448 ;
        RECT 0.27 0.178 0.515 0.1967 ;
        RECT 0.338 0.1227 0.626 0.1413 ;
        RECT 0.626 0.1227 0.654 0.1413 ;
        RECT 0.626 0.1413 0.654 0.184 ;
        RECT 0.392 0.424 0.754 0.4453 ;
        RECT 0.754 0.1647 0.782 0.364 ;
        RECT 0.466 0.0679 0.878 0.0867 ;
        RECT 1.061 0.16 1.098 0.2973 ;
        RECT 1.202 0.114 1.23 0.3407 ;
        RECT 1.458 0.0973 1.49 0.4653 ;
        RECT 1.165 0.412 1.33 0.4307 ;
        RECT 1.33 0.0427 1.358 0.0613 ;
        RECT 1.33 0.0613 1.358 0.244 ;
        RECT 1.33 0.244 1.358 0.412 ;
        RECT 1.33 0.412 1.358 0.4307 ;
        RECT 1.358 0.0427 1.607 0.0613 ;
        RECT 1.607 0.0427 1.635 0.0613 ;
        RECT 1.607 0.0613 1.635 0.244 ;
        RECT 1.554 0.3067 1.582 0.416 ;
        RECT 1.554 0.416 1.582 0.4533 ;
        RECT 1.582 0.416 1.714 0.4533 ;
        RECT 1.714 0.048 1.742 0.3067 ;
        RECT 1.714 0.3067 1.742 0.416 ;
        RECT 1.714 0.416 1.742 0.4533 ;
        RECT 0.178 0.0833 0.206 0.3827 ;
        RECT 0.6899 0.258 0.718 0.3933 ;
        RECT 0.8179 0.1713 0.85 0.3127 ;
        RECT 0.6899 0.1107 0.718 0.1293 ;
        RECT 0.6899 0.1293 0.718 0.184 ;
        RECT 0.718 0.1107 0.942 0.1293 ;
        RECT 0.991 0.1613 1.025 0.2813 ;
        RECT 0.79 0.424 1.066 0.4453 ;
        RECT 0.904 0.1827 0.932 0.3267 ;
        RECT 0.904 0.3267 0.932 0.3453 ;
        RECT 0.932 0.3267 1.1339 0.3453 ;
        RECT 1.1339 0.0547 1.166 0.1827 ;
        RECT 1.1339 0.1827 1.166 0.3267 ;
        RECT 1.1339 0.3267 1.166 0.3453 ;
        RECT 1.266 0.1187 1.294 0.3827 ;
        RECT 1.3939 0.1187 1.422 0.3293 ;
        RECT 1.532 0.1027 1.571 0.2773 ;
      LAYER V1 ;
        RECT 0.114 0.1827 0.1419 0.2013 ;
        RECT 0.178 0.3533 0.206 0.372 ;
        RECT 0.6899 0.3533 0.718 0.372 ;
        RECT 0.754 0.268 0.782 0.2867 ;
        RECT 0.8179 0.1827 0.846 0.2013 ;
        RECT 0.997 0.2253 1.025 0.244 ;
        RECT 1.061 0.268 1.089 0.2867 ;
        RECT 1.202 0.1827 1.23 0.2013 ;
        RECT 1.266 0.3533 1.294 0.372 ;
        RECT 1.3939 0.1827 1.422 0.2013 ;
        RECT 1.532 0.2253 1.56 0.244 ;
      LAYER M1 ;
        RECT 0.045 0.064 0.083 0.1359 ;
        RECT 0.045 0.1359 0.083 0.1547 ;
        RECT 0.045 0.4027 0.083 0.4213 ;
        RECT 0.045 0.4213 0.083 0.4586 ;
        RECT 0.083 0.1359 0.114 0.1547 ;
        RECT 0.083 0.4027 0.114 0.4213 ;
        RECT 0.114 0.1359 0.1419 0.1547 ;
        RECT 0.114 0.1547 0.1419 0.4027 ;
        RECT 0.114 0.4027 0.1419 0.4213 ;
        RECT 0.242 0.064 0.27 0.178 ;
        RECT 0.242 0.178 0.27 0.1967 ;
        RECT 0.242 0.1967 0.27 0.448 ;
        RECT 0.27 0.178 0.515 0.1967 ;
        RECT 0.338 0.1227 0.626 0.1413 ;
        RECT 0.626 0.1227 0.654 0.1413 ;
        RECT 0.626 0.1413 0.654 0.184 ;
        RECT 0.392 0.424 0.754 0.4453 ;
        RECT 0.754 0.1647 0.782 0.364 ;
        RECT 0.466 0.0679 0.878 0.0867 ;
        RECT 1.061 0.16 1.098 0.2973 ;
        RECT 1.202 0.114 1.23 0.3407 ;
        RECT 1.458 0.0973 1.49 0.4653 ;
        RECT 1.165 0.412 1.33 0.4307 ;
        RECT 1.33 0.0427 1.358 0.0613 ;
        RECT 1.33 0.0613 1.358 0.244 ;
        RECT 1.33 0.244 1.358 0.412 ;
        RECT 1.33 0.412 1.358 0.4307 ;
        RECT 1.358 0.0427 1.607 0.0613 ;
        RECT 1.607 0.0427 1.635 0.0613 ;
        RECT 1.607 0.0613 1.635 0.244 ;
        RECT 1.554 0.3067 1.582 0.416 ;
        RECT 1.554 0.416 1.582 0.4533 ;
        RECT 1.582 0.416 1.714 0.4533 ;
        RECT 1.714 0.048 1.742 0.3067 ;
        RECT 1.714 0.3067 1.742 0.416 ;
        RECT 1.714 0.416 1.742 0.4533 ;
        RECT 0.178 0.0833 0.206 0.3827 ;
        RECT 0.6899 0.258 0.718 0.3933 ;
        RECT 0.8179 0.1713 0.85 0.3127 ;
        RECT 0.6899 0.1107 0.718 0.1293 ;
        RECT 0.6899 0.1293 0.718 0.184 ;
        RECT 0.718 0.1107 0.942 0.1293 ;
        RECT 0.991 0.1613 1.025 0.2813 ;
        RECT 0.79 0.424 1.066 0.4453 ;
        RECT 0.904 0.1827 0.932 0.3267 ;
        RECT 0.904 0.3267 0.932 0.3453 ;
        RECT 0.932 0.3267 1.1339 0.3453 ;
        RECT 1.1339 0.0547 1.166 0.1827 ;
        RECT 1.1339 0.1827 1.166 0.3267 ;
        RECT 1.1339 0.3267 1.166 0.3453 ;
        RECT 1.266 0.1187 1.294 0.3827 ;
        RECT 1.3939 0.1187 1.422 0.3293 ;
        RECT 1.532 0.1027 1.571 0.2773 ;
  END
END SDFFRNQ_X1_8T

MACRO SDFFSNQ_X1_8T
  CLASS core ;
  FOREIGN SDFFSNQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.92 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.256 0.51 0.352 ;
        RECT 0.51 0.256 0.526 0.352 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.248 0.334 0.3813 ;
        RECT 0.306 0.3813 0.334 0.4 ;
        RECT 0.334 0.3813 0.51 0.4 ;
        RECT 0.51 0.3813 0.562 0.4 ;
        RECT 0.562 0.2093 0.59 0.248 ;
        RECT 0.562 0.248 0.59 0.3813 ;
        RECT 0.562 0.3813 0.59 0.4 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.242 0.398 0.3413 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.958 0.2253 1.454 0.244 ;
        RECT 1.454 0.2253 1.586 0.244 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1813 0.078 0.3413 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.0427 1.872 0.4693 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.49336 0.5307 ;
        RECT 0.49336 0.4933 0.782 0.5307 ;
        RECT 0.782 0.4933 0.862 0.5307 ;
        RECT 0.862 0.4933 1.646 0.5307 ;
        RECT 1.646 0.4933 1.742 0.5307 ;
        RECT 1.742 0.4933 1.93 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.93 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.3533 1.326 0.372 ;
        RECT 0.722 0.268 1.114 0.2867 ;
        RECT 0.082 0.1827 1.454 0.2013 ;
      LAYER MINT1 ;
        RECT 0.146 0.3533 1.326 0.372 ;
        RECT 0.722 0.268 1.114 0.2867 ;
        RECT 0.082 0.1827 1.454 0.2013 ;
      LAYER M1 ;
        RECT 0.048 0.0427 0.08 0.1333 ;
        RECT 0.048 0.1333 0.08 0.133328 ;
        RECT 0.048 0.4027 0.08 0.4213 ;
        RECT 0.048 0.4213 0.08 0.4586 ;
        RECT 0.08 0.1333 0.114 0.133328 ;
        RECT 0.08 0.4027 0.114 0.4213 ;
        RECT 0.114 0.1333 0.1419 0.133328 ;
        RECT 0.114 0.152 0.1419 0.4027 ;
        RECT 0.114 0.4027 0.1419 0.4213 ;
        RECT 0.242 0.0547 0.27 0.1773 ;
        RECT 0.242 0.1773 0.27 0.1967 ;
        RECT 0.242 0.1967 0.27 0.1973 ;
        RECT 0.242 0.1973 0.27 0.4573 ;
        RECT 0.27 0.1773 0.434 0.1967 ;
        RECT 0.434 0.1773 0.51 0.1967 ;
        RECT 0.434 0.1967 0.51 0.1973 ;
        RECT 0.338 0.1227 0.626 0.1413 ;
        RECT 0.626 0.1227 0.654 0.1413 ;
        RECT 0.626 0.1413 0.654 0.184 ;
        RECT 0.392 0.424 0.746 0.4453 ;
        RECT 0.754 0.1587 0.782 0.3647 ;
        RECT 0.466 0.0679 0.878 0.0867 ;
        RECT 0.98 0.2147 1.018 0.2793 ;
        RECT 0.898 0.1827 0.926 0.3247 ;
        RECT 0.898 0.3247 0.926 0.3433 ;
        RECT 0.926 0.3247 1.008 0.3433 ;
        RECT 1.008 0.3247 1.04 0.3433 ;
        RECT 1.008 0.3433 1.04 0.4693 ;
        RECT 1.04 0.3247 1.1379 0.3433 ;
        RECT 1.1379 0.0653 1.166 0.1827 ;
        RECT 1.1379 0.1827 1.166 0.3247 ;
        RECT 1.1379 0.3247 1.166 0.3433 ;
        RECT 1.266 0.1187 1.294 0.3827 ;
        RECT 1.3939 0.1187 1.422 0.268 ;
        RECT 1.526 0.1227 1.554 0.2687 ;
        RECT 1.402 0.4253 1.646 0.444 ;
        RECT 0.178 0.064 0.206 0.4127 ;
        RECT 0.654 0.258 0.682 0.3827 ;
        RECT 0.83 0.1713 0.862 0.3127 ;
        RECT 0.6899 0.1107 0.718 0.1293 ;
        RECT 0.6899 0.1293 0.718 0.184 ;
        RECT 0.718 0.1107 0.942 0.1293 ;
        RECT 1.054 0.16 1.092 0.2973 ;
        RECT 1.202 0.114 1.23 0.2553 ;
        RECT 1.165 0.412 1.33 0.4307 ;
        RECT 1.33 0.0547 1.358 0.0733 ;
        RECT 1.33 0.0733 1.358 0.244 ;
        RECT 1.33 0.244 1.358 0.412 ;
        RECT 1.33 0.412 1.358 0.4307 ;
        RECT 1.358 0.0547 1.607 0.0733 ;
        RECT 1.607 0.0547 1.645 0.0733 ;
        RECT 1.607 0.0733 1.645 0.244 ;
        RECT 1.462 0.268 1.49 0.3827 ;
        RECT 1.462 0.3827 1.49 0.4013 ;
        RECT 1.49 0.3827 1.714 0.4013 ;
        RECT 1.714 0.064 1.742 0.268 ;
        RECT 1.714 0.268 1.742 0.3827 ;
        RECT 1.714 0.3827 1.742 0.4013 ;
      LAYER V1 ;
        RECT 0.114 0.1827 0.1419 0.2013 ;
        RECT 0.178 0.3533 0.206 0.372 ;
        RECT 0.654 0.3533 0.682 0.372 ;
        RECT 0.754 0.268 0.782 0.2867 ;
        RECT 0.834 0.1827 0.862 0.2013 ;
        RECT 0.99 0.2253 1.018 0.244 ;
        RECT 1.054 0.268 1.082 0.2867 ;
        RECT 1.202 0.1827 1.23 0.2013 ;
        RECT 1.266 0.3533 1.294 0.372 ;
        RECT 1.3939 0.1827 1.422 0.2013 ;
        RECT 1.526 0.2253 1.554 0.244 ;
      LAYER M1 ;
        RECT 0.048 0.0427 0.08 0.1333 ;
        RECT 0.048 0.1333 0.08 0.133328 ;
        RECT 0.048 0.4027 0.08 0.4213 ;
        RECT 0.048 0.4213 0.08 0.4586 ;
        RECT 0.08 0.1333 0.114 0.133328 ;
        RECT 0.08 0.4027 0.114 0.4213 ;
        RECT 0.114 0.1333 0.1419 0.133328 ;
        RECT 0.114 0.152 0.1419 0.4027 ;
        RECT 0.114 0.4027 0.1419 0.4213 ;
        RECT 0.242 0.0547 0.27 0.1773 ;
        RECT 0.242 0.1773 0.27 0.1967 ;
        RECT 0.242 0.1967 0.27 0.1973 ;
        RECT 0.242 0.1973 0.27 0.4573 ;
        RECT 0.27 0.1773 0.434 0.1967 ;
        RECT 0.434 0.1773 0.51 0.1967 ;
        RECT 0.434 0.1967 0.51 0.1973 ;
        RECT 0.338 0.1227 0.626 0.1413 ;
        RECT 0.626 0.1227 0.654 0.1413 ;
        RECT 0.626 0.1413 0.654 0.184 ;
        RECT 0.392 0.424 0.746 0.4453 ;
        RECT 0.754 0.1587 0.782 0.3647 ;
        RECT 0.466 0.0679 0.878 0.0867 ;
        RECT 0.98 0.2147 1.018 0.2793 ;
        RECT 0.898 0.1827 0.926 0.3247 ;
        RECT 0.898 0.3247 0.926 0.3433 ;
        RECT 0.926 0.3247 1.008 0.3433 ;
        RECT 1.008 0.3247 1.04 0.3433 ;
        RECT 1.008 0.3433 1.04 0.4693 ;
        RECT 1.04 0.3247 1.1379 0.3433 ;
        RECT 1.1379 0.0653 1.166 0.1827 ;
        RECT 1.1379 0.1827 1.166 0.3247 ;
        RECT 1.1379 0.3247 1.166 0.3433 ;
        RECT 1.266 0.1187 1.294 0.3827 ;
        RECT 1.3939 0.1187 1.422 0.268 ;
        RECT 1.526 0.1227 1.554 0.2687 ;
        RECT 1.402 0.4253 1.646 0.444 ;
        RECT 0.178 0.064 0.206 0.4127 ;
        RECT 0.654 0.258 0.682 0.3827 ;
        RECT 0.83 0.1713 0.862 0.3127 ;
        RECT 0.6899 0.1107 0.718 0.1293 ;
        RECT 0.6899 0.1293 0.718 0.184 ;
        RECT 0.718 0.1107 0.942 0.1293 ;
        RECT 1.054 0.16 1.092 0.2973 ;
        RECT 1.202 0.114 1.23 0.2553 ;
        RECT 1.165 0.412 1.33 0.4307 ;
        RECT 1.33 0.0547 1.358 0.0733 ;
        RECT 1.33 0.0733 1.358 0.244 ;
        RECT 1.33 0.244 1.358 0.412 ;
        RECT 1.33 0.412 1.358 0.4307 ;
        RECT 1.358 0.0547 1.607 0.0733 ;
        RECT 1.607 0.0547 1.645 0.0733 ;
        RECT 1.607 0.0733 1.645 0.244 ;
        RECT 1.462 0.268 1.49 0.3827 ;
        RECT 1.462 0.3827 1.49 0.4013 ;
        RECT 1.49 0.3827 1.714 0.4013 ;
        RECT 1.714 0.064 1.742 0.268 ;
        RECT 1.714 0.268 1.742 0.3827 ;
        RECT 1.714 0.3827 1.742 0.4013 ;
  END
END SDFFSNQ_X1_8T

MACRO TBUF_X1_8T
  CLASS core ;
  FOREIGN TBUF_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.328 ;
        RECT 0.114 0.328 0.1419 0.3467 ;
        RECT 0.1419 0.328 0.206 0.3467 ;
        RECT 0.206 0.328 0.242 0.3467 ;
        RECT 0.242 0.204 0.27 0.256 ;
        RECT 0.242 0.256 0.27 0.328 ;
        RECT 0.242 0.328 0.27 0.3467 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.2467 0.462 0.384 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.0427 0.656 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.588 0.5307 ;
        RECT 0.588 0.4933 0.714 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.714 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2787 ;
        RECT 0.05 0.2787 0.078 0.4573 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2787 ;
        RECT 0.146 0.3827 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3827 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3827 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.2093 ;
        RECT 0.306 0.2093 0.334 0.3827 ;
        RECT 0.306 0.3827 0.334 0.4013 ;
        RECT 0.334 0.0679 0.51 0.0867 ;
        RECT 0.51 0.0679 0.542 0.0867 ;
        RECT 0.51 0.0867 0.542 0.1533 ;
        RECT 0.51 0.1533 0.542 0.172 ;
        RECT 0.51 0.172 0.542 0.2093 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2507 ;
        RECT 0.37 0.2507 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.56 0.444 ;
        RECT 0.56 0.2507 0.588 0.4253 ;
        RECT 0.56 0.4253 0.588 0.444 ;
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2787 ;
        RECT 0.05 0.2787 0.078 0.4573 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2787 ;
        RECT 0.146 0.3827 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3827 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3827 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.2093 ;
        RECT 0.306 0.2093 0.334 0.3827 ;
        RECT 0.306 0.3827 0.334 0.4013 ;
        RECT 0.334 0.0679 0.51 0.0867 ;
        RECT 0.51 0.0679 0.542 0.0867 ;
        RECT 0.51 0.0867 0.542 0.1533 ;
        RECT 0.51 0.1533 0.542 0.172 ;
        RECT 0.51 0.172 0.542 0.2093 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2507 ;
        RECT 0.37 0.2507 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.56 0.444 ;
        RECT 0.56 0.2507 0.588 0.4253 ;
        RECT 0.56 0.4253 0.588 0.444 ;
  END
END TBUF_X1_8T

MACRO TBUF_X2_8T
  CLASS core ;
  FOREIGN TBUF_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.336 ;
        RECT 0.114 0.336 0.1419 0.3547 ;
        RECT 0.1419 0.336 0.206 0.3547 ;
        RECT 0.206 0.336 0.242 0.3547 ;
        RECT 0.242 0.204 0.27 0.256 ;
        RECT 0.242 0.256 0.27 0.336 ;
        RECT 0.242 0.336 0.27 0.3547 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.2547 0.462 0.384 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.0467 0.656 0.4639 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.53 0.5307 ;
        RECT 0.53 0.4933 0.778 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.778 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.408 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.146 0.3786 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3786 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3786 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.2093 ;
        RECT 0.306 0.2093 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4013 ;
        RECT 0.334 0.0679 0.482 0.0867 ;
        RECT 0.482 0.0679 0.514 0.0867 ;
        RECT 0.482 0.0867 0.514 0.1533 ;
        RECT 0.482 0.1533 0.514 0.172 ;
        RECT 0.482 0.172 0.514 0.2093 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2953 ;
        RECT 0.37 0.2953 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.498 0.444 ;
        RECT 0.498 0.2953 0.53 0.4253 ;
        RECT 0.498 0.4253 0.53 0.444 ;
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.408 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.146 0.3786 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3786 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3786 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.2093 ;
        RECT 0.306 0.2093 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4013 ;
        RECT 0.334 0.0679 0.482 0.0867 ;
        RECT 0.482 0.0679 0.514 0.0867 ;
        RECT 0.482 0.0867 0.514 0.1533 ;
        RECT 0.482 0.1533 0.514 0.172 ;
        RECT 0.482 0.172 0.514 0.2093 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2953 ;
        RECT 0.37 0.2953 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.498 0.444 ;
        RECT 0.498 0.2953 0.53 0.4253 ;
        RECT 0.498 0.4253 0.53 0.444 ;
  END
END TBUF_X2_8T

MACRO TBUF_X4_8T
  CLASS core ;
  FOREIGN TBUF_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.96 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.3227 ;
        RECT 0.114 0.3227 0.1419 0.3413 ;
        RECT 0.1419 0.3227 0.206 0.3413 ;
        RECT 0.206 0.3227 0.242 0.3413 ;
        RECT 0.242 0.204 0.27 0.256 ;
        RECT 0.242 0.256 0.27 0.3227 ;
        RECT 0.242 0.3227 0.27 0.3413 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.2306 0.462 0.396 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.6879 0.0427 0.72 0.1493 ;
        RECT 0.6879 0.1493 0.72 0.1707 ;
        RECT 0.6879 0.3413 0.72 0.36 ;
        RECT 0.6879 0.36 0.72 0.3806 ;
        RECT 0.6879 0.3806 0.72 0.4693 ;
        RECT 0.72 0.1493 0.8129 0.1707 ;
        RECT 0.72 0.3413 0.8129 0.36 ;
        RECT 0.8129 0.0427 0.8139 0.1493 ;
        RECT 0.8129 0.1493 0.8139 0.1707 ;
        RECT 0.8129 0.3413 0.8139 0.36 ;
        RECT 0.8139 0.0427 0.8159 0.1493 ;
        RECT 0.8139 0.1493 0.8159 0.1707 ;
        RECT 0.8139 0.3413 0.8159 0.36 ;
        RECT 0.8159 0.0427 0.838 0.1493 ;
        RECT 0.8159 0.1493 0.838 0.1707 ;
        RECT 0.8159 0.3413 0.838 0.36 ;
        RECT 0.8159 0.36 0.838 0.3806 ;
        RECT 0.8159 0.3806 0.838 0.4693 ;
        RECT 0.838 0.0427 0.848 0.1493 ;
        RECT 0.838 0.1493 0.848 0.1707 ;
        RECT 0.838 0.3413 0.848 0.36 ;
        RECT 0.838 0.36 0.848 0.3806 ;
        RECT 0.838 0.3806 0.848 0.4693 ;
        RECT 0.848 0.0427 0.851 0.1493 ;
        RECT 0.848 0.1493 0.851 0.1707 ;
        RECT 0.848 0.3413 0.851 0.36 ;
        RECT 0.848 0.36 0.851 0.3806 ;
        RECT 0.851 0.1493 0.882 0.1707 ;
        RECT 0.851 0.3413 0.882 0.36 ;
        RECT 0.851 0.36 0.882 0.3806 ;
        RECT 0.882 0.1493 0.91 0.1707 ;
        RECT 0.882 0.1707 0.91 0.3413 ;
        RECT 0.882 0.3413 0.91 0.36 ;
        RECT 0.882 0.36 0.91 0.3806 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.8139 0.5307 ;
        RECT 0.8139 0.4933 0.838 0.5307 ;
        RECT 0.838 0.4933 0.97 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.97 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2587 ;
        RECT 0.37 0.2587 0.398 0.276 ;
        RECT 0.37 0.276 0.398 0.3053 ;
        RECT 0.37 0.3053 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.526 0.444 ;
        RECT 0.526 0.2587 0.582 0.276 ;
        RECT 0.526 0.276 0.582 0.3053 ;
        RECT 0.526 0.3053 0.582 0.4253 ;
        RECT 0.526 0.4253 0.582 0.444 ;
        RECT 0.582 0.276 0.8139 0.3053 ;
        RECT 0.05 0.064 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.396 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.146 0.3786 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3786 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3786 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.1947 ;
        RECT 0.306 0.1947 0.334 0.2133 ;
        RECT 0.306 0.2133 0.334 0.2347 ;
        RECT 0.306 0.2347 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4013 ;
        RECT 0.334 0.0679 0.526 0.0867 ;
        RECT 0.526 0.0679 0.582 0.0867 ;
        RECT 0.526 0.0867 0.582 0.1533 ;
        RECT 0.526 0.1533 0.582 0.172 ;
        RECT 0.526 0.172 0.582 0.1947 ;
        RECT 0.526 0.1947 0.582 0.2133 ;
        RECT 0.526 0.2133 0.582 0.2347 ;
        RECT 0.582 0.1947 0.838 0.2133 ;
      LAYER M1 ;
        RECT 0.082 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2587 ;
        RECT 0.37 0.2587 0.398 0.276 ;
        RECT 0.37 0.276 0.398 0.3053 ;
        RECT 0.37 0.3053 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.526 0.444 ;
        RECT 0.526 0.2587 0.582 0.276 ;
        RECT 0.526 0.276 0.582 0.3053 ;
        RECT 0.526 0.3053 0.582 0.4253 ;
        RECT 0.526 0.4253 0.582 0.444 ;
        RECT 0.582 0.276 0.8139 0.3053 ;
        RECT 0.05 0.064 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.396 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.146 0.3786 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3786 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3786 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.1947 ;
        RECT 0.306 0.1947 0.334 0.2133 ;
        RECT 0.306 0.2133 0.334 0.2347 ;
        RECT 0.306 0.2347 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4013 ;
        RECT 0.334 0.0679 0.526 0.0867 ;
        RECT 0.526 0.0679 0.582 0.0867 ;
        RECT 0.526 0.0867 0.582 0.1533 ;
        RECT 0.526 0.1533 0.582 0.172 ;
        RECT 0.526 0.172 0.582 0.1947 ;
        RECT 0.526 0.1947 0.582 0.2133 ;
        RECT 0.526 0.2133 0.582 0.2347 ;
        RECT 0.582 0.1947 0.838 0.2133 ;
  END
END TBUF_X4_8T

MACRO TBUF_X8_8T
  CLASS core ;
  FOREIGN TBUF_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.344 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.3227 ;
        RECT 0.114 0.3227 0.1419 0.3413 ;
        RECT 0.1419 0.3227 0.222 0.3413 ;
        RECT 0.222 0.3227 0.306 0.3413 ;
        RECT 0.306 0.2133 0.334 0.256 ;
        RECT 0.306 0.256 0.334 0.3227 ;
        RECT 0.306 0.3227 0.334 0.3413 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.2306 0.526 0.268 ;
        RECT 0.498 0.268 0.526 0.2893 ;
        RECT 0.498 0.2893 0.526 0.384 ;
        RECT 0.526 0.268 0.622 0.2893 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8159 0.0427 0.848 0.0887 ;
        RECT 0.8159 0.0887 0.848 0.1067 ;
        RECT 0.8159 0.1067 0.848 0.128 ;
        RECT 0.8159 0.346 0.848 0.3847 ;
        RECT 0.8159 0.3847 0.848 0.3853 ;
        RECT 0.8159 0.3853 0.848 0.4693 ;
        RECT 0.848 0.1067 1.183 0.128 ;
        RECT 0.848 0.346 1.183 0.3847 ;
        RECT 1.183 0.1067 1.198 0.128 ;
        RECT 1.183 0.346 1.198 0.3847 ;
        RECT 1.198 0.1067 1.2 0.128 ;
        RECT 1.198 0.346 1.2 0.3847 ;
        RECT 1.2 0.0427 1.232 0.0887 ;
        RECT 1.2 0.0887 1.232 0.1067 ;
        RECT 1.2 0.1067 1.232 0.128 ;
        RECT 1.2 0.346 1.232 0.3847 ;
        RECT 1.2 0.3847 1.232 0.3853 ;
        RECT 1.2 0.3853 1.232 0.4693 ;
        RECT 1.232 0.0887 1.266 0.1067 ;
        RECT 1.232 0.1067 1.266 0.128 ;
        RECT 1.232 0.346 1.266 0.3847 ;
        RECT 1.232 0.3847 1.266 0.3853 ;
        RECT 1.266 0.0887 1.294 0.1067 ;
        RECT 1.266 0.1067 1.294 0.128 ;
        RECT 1.266 0.128 1.294 0.346 ;
        RECT 1.266 0.346 1.294 0.3847 ;
        RECT 1.266 0.3847 1.294 0.3853 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.183 0.5307 ;
        RECT 1.183 0.4933 1.198 0.5307 ;
        RECT 1.198 0.4933 1.354 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.354 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2867 ;
        RECT 0.05 0.2867 0.078 0.4253 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.222 0.2267 ;
        RECT 0.178 0.2267 0.222 0.2867 ;
        RECT 0.146 0.3827 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3827 0.23 0.4013 ;
        RECT 0.23 0.0679 0.37 0.0867 ;
        RECT 0.1533 0.1533 0.37 0.172 ;
        RECT 0.23 0.3827 0.37 0.4013 ;
        RECT 0.37 0.0679 0.398 0.0867 ;
        RECT 0.37 0.1533 0.398 0.172 ;
        RECT 0.37 0.172 0.398 0.1906 ;
        RECT 0.37 0.1906 0.398 0.228 ;
        RECT 0.37 0.228 0.398 0.3827 ;
        RECT 0.37 0.3827 0.398 0.4013 ;
        RECT 0.398 0.0679 0.6899 0.0867 ;
        RECT 0.6899 0.0679 0.718 0.0867 ;
        RECT 0.6899 0.0867 0.718 0.1533 ;
        RECT 0.6899 0.1533 0.718 0.172 ;
        RECT 0.6899 0.172 0.718 0.1906 ;
        RECT 0.6899 0.1906 0.718 0.228 ;
        RECT 0.718 0.172 1.198 0.1906 ;
        RECT 0.122 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.434 0.1293 ;
        RECT 0.274 0.4253 0.434 0.444 ;
        RECT 0.434 0.1107 0.462 0.1293 ;
        RECT 0.434 0.1293 0.462 0.2573 ;
        RECT 0.434 0.2573 0.462 0.2687 ;
        RECT 0.434 0.2687 0.462 0.3073 ;
        RECT 0.434 0.3073 0.462 0.4253 ;
        RECT 0.434 0.4253 0.462 0.444 ;
        RECT 0.462 0.4253 0.66 0.444 ;
        RECT 0.66 0.2573 0.718 0.2687 ;
        RECT 0.66 0.2687 0.718 0.3073 ;
        RECT 0.66 0.3073 0.718 0.4253 ;
        RECT 0.66 0.4253 0.718 0.444 ;
        RECT 0.718 0.2687 1.183 0.3073 ;
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2867 ;
        RECT 0.05 0.2867 0.078 0.4253 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.222 0.2267 ;
        RECT 0.178 0.2267 0.222 0.2867 ;
        RECT 0.146 0.3827 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3827 0.23 0.4013 ;
        RECT 0.23 0.0679 0.37 0.0867 ;
        RECT 0.1533 0.1533 0.37 0.172 ;
        RECT 0.23 0.3827 0.37 0.4013 ;
        RECT 0.37 0.0679 0.398 0.0867 ;
        RECT 0.37 0.1533 0.398 0.172 ;
        RECT 0.37 0.172 0.398 0.1906 ;
        RECT 0.37 0.1906 0.398 0.228 ;
        RECT 0.37 0.228 0.398 0.3827 ;
        RECT 0.37 0.3827 0.398 0.4013 ;
        RECT 0.398 0.0679 0.6899 0.0867 ;
        RECT 0.6899 0.0679 0.718 0.0867 ;
        RECT 0.6899 0.0867 0.718 0.1533 ;
        RECT 0.6899 0.1533 0.718 0.172 ;
        RECT 0.6899 0.172 0.718 0.1906 ;
        RECT 0.6899 0.1906 0.718 0.228 ;
        RECT 0.718 0.172 1.198 0.1906 ;
        RECT 0.122 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.434 0.1293 ;
        RECT 0.274 0.4253 0.434 0.444 ;
        RECT 0.434 0.1107 0.462 0.1293 ;
        RECT 0.434 0.1293 0.462 0.2573 ;
        RECT 0.434 0.2573 0.462 0.2687 ;
        RECT 0.434 0.2687 0.462 0.3073 ;
        RECT 0.434 0.3073 0.462 0.4253 ;
        RECT 0.434 0.4253 0.462 0.444 ;
        RECT 0.462 0.4253 0.66 0.444 ;
        RECT 0.66 0.2573 0.718 0.2687 ;
        RECT 0.66 0.2687 0.718 0.3073 ;
        RECT 0.66 0.3073 0.718 0.4253 ;
        RECT 0.66 0.4253 0.718 0.444 ;
        RECT 0.718 0.2687 1.183 0.3073 ;
  END
END TBUF_X8_8T

MACRO TBUF_X12_8T
  CLASS core ;
  FOREIGN TBUF_X12_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.728 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.34 ;
        RECT 0.114 0.34 0.1419 0.3587 ;
        RECT 0.1419 0.34 0.206 0.3587 ;
        RECT 0.206 0.34 0.242 0.3587 ;
        RECT 0.242 0.204 0.27 0.256 ;
        RECT 0.242 0.256 0.27 0.34 ;
        RECT 0.242 0.34 0.27 0.3587 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.268 0.498 0.2987 ;
        RECT 0.498 0.2306 0.526 0.268 ;
        RECT 0.498 0.268 0.526 0.2987 ;
        RECT 0.526 0.268 0.626 0.2987 ;
        RECT 0.626 0.268 0.654 0.2987 ;
        RECT 0.626 0.2987 0.654 0.384 ;
        RECT 0.654 0.268 0.71 0.2987 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.684 0.5307 ;
        RECT 1.684 0.4933 1.738 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.738 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2373 ;
        RECT 0.37 0.2373 0.398 0.252 ;
        RECT 0.37 0.252 0.398 0.284 ;
        RECT 0.37 0.284 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.783 0.444 ;
        RECT 0.783 0.2373 0.839 0.252 ;
        RECT 0.783 0.252 0.839 0.284 ;
        RECT 0.783 0.284 0.839 0.4253 ;
        RECT 0.783 0.4253 0.839 0.444 ;
        RECT 0.839 0.252 1.557 0.284 ;
        RECT 0.882 0.0679 0.931 0.0867 ;
        RECT 0.931 0.0679 0.989 0.0867 ;
        RECT 0.931 0.3547 0.989 0.3759 ;
        RECT 0.931 0.3759 0.989 0.4133 ;
        RECT 0.989 0.0679 1.572 0.0867 ;
        RECT 0.989 0.3547 1.572 0.3759 ;
        RECT 1.572 0.0487 1.586 0.0679 ;
        RECT 1.572 0.0679 1.586 0.0867 ;
        RECT 1.572 0.3547 1.586 0.3759 ;
        RECT 1.586 0.0487 1.614 0.0679 ;
        RECT 1.586 0.0679 1.614 0.0867 ;
        RECT 1.586 0.3547 1.614 0.3759 ;
        RECT 1.586 0.3759 1.614 0.4133 ;
        RECT 1.586 0.4133 1.614 0.41334 ;
        RECT 1.614 0.0487 1.6279 0.0679 ;
        RECT 1.614 0.0679 1.6279 0.0867 ;
        RECT 1.614 0.3547 1.6279 0.3759 ;
        RECT 1.6279 0.0679 1.629 0.0867 ;
        RECT 1.6279 0.3547 1.629 0.3759 ;
        RECT 1.629 0.0679 1.684 0.0867 ;
        RECT 1.629 0.0867 1.684 0.3547 ;
        RECT 1.629 0.3547 1.684 0.3759 ;
        RECT 0.05 0.1159 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.448 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.1419 0.0679 0.146 0.0867 ;
        RECT 0.1419 0.0867 0.146 0.1533 ;
        RECT 0.1419 0.1533 0.146 0.1667 ;
        RECT 0.1419 0.1667 0.146 0.16678 ;
        RECT 0.146 0.0679 0.17 0.0867 ;
        RECT 0.146 0.0867 0.17 0.1533 ;
        RECT 0.146 0.1533 0.17 0.1667 ;
        RECT 0.146 0.1667 0.17 0.16678 ;
        RECT 0.146 0.3827 0.17 0.4013 ;
        RECT 0.17 0.0679 0.306 0.0867 ;
        RECT 0.17 0.1533 0.306 0.1667 ;
        RECT 0.17 0.1667 0.306 0.16678 ;
        RECT 0.17 0.3827 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.1667 ;
        RECT 0.306 0.1667 0.334 0.16678 ;
        RECT 0.306 0.172 0.334 0.196 ;
        RECT 0.306 0.196 0.334 0.3827 ;
        RECT 0.306 0.3827 0.334 0.4013 ;
        RECT 0.334 0.0679 0.782 0.0867 ;
        RECT 0.782 0.0679 0.8139 0.0867 ;
        RECT 0.782 0.0867 0.8139 0.1533 ;
        RECT 0.782 0.1533 0.8139 0.1667 ;
        RECT 0.782 0.1667 0.8139 0.16678 ;
        RECT 0.782 0.172 0.8139 0.196 ;
        RECT 0.8139 0.1667 1.593 0.16678 ;
        RECT 0.8139 0.172 1.593 0.196 ;
      LAYER M1 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2373 ;
        RECT 0.37 0.2373 0.398 0.252 ;
        RECT 0.37 0.252 0.398 0.284 ;
        RECT 0.37 0.284 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.783 0.444 ;
        RECT 0.783 0.2373 0.839 0.252 ;
        RECT 0.783 0.252 0.839 0.284 ;
        RECT 0.783 0.284 0.839 0.4253 ;
        RECT 0.783 0.4253 0.839 0.444 ;
        RECT 0.839 0.252 1.557 0.284 ;
        RECT 0.882 0.0679 0.931 0.0867 ;
        RECT 0.931 0.0679 0.989 0.0867 ;
        RECT 0.931 0.3547 0.989 0.3759 ;
        RECT 0.931 0.3759 0.989 0.4133 ;
        RECT 0.989 0.0679 1.572 0.0867 ;
        RECT 0.989 0.3547 1.572 0.3759 ;
        RECT 1.572 0.0487 1.586 0.0679 ;
        RECT 1.572 0.0679 1.586 0.0867 ;
        RECT 1.572 0.3547 1.586 0.3759 ;
        RECT 1.586 0.0487 1.614 0.0679 ;
        RECT 1.586 0.0679 1.614 0.0867 ;
        RECT 1.586 0.3547 1.614 0.3759 ;
        RECT 1.586 0.3759 1.614 0.4133 ;
        RECT 1.586 0.4133 1.614 0.41334 ;
        RECT 1.614 0.0487 1.6279 0.0679 ;
        RECT 1.614 0.0679 1.6279 0.0867 ;
        RECT 1.614 0.3547 1.6279 0.3759 ;
        RECT 1.6279 0.0679 1.629 0.0867 ;
        RECT 1.6279 0.3547 1.629 0.3759 ;
        RECT 1.629 0.0679 1.684 0.0867 ;
        RECT 1.629 0.0867 1.684 0.3547 ;
        RECT 1.629 0.3547 1.684 0.3759 ;
        RECT 0.05 0.1159 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.448 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.1419 0.0679 0.146 0.0867 ;
        RECT 0.1419 0.0867 0.146 0.1533 ;
        RECT 0.1419 0.1533 0.146 0.1667 ;
        RECT 0.1419 0.1667 0.146 0.16678 ;
        RECT 0.146 0.0679 0.17 0.0867 ;
        RECT 0.146 0.0867 0.17 0.1533 ;
        RECT 0.146 0.1533 0.17 0.1667 ;
        RECT 0.146 0.1667 0.17 0.16678 ;
        RECT 0.146 0.3827 0.17 0.4013 ;
        RECT 0.17 0.0679 0.306 0.0867 ;
        RECT 0.17 0.1533 0.306 0.1667 ;
        RECT 0.17 0.1667 0.306 0.16678 ;
        RECT 0.17 0.3827 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.1667 ;
        RECT 0.306 0.1667 0.334 0.16678 ;
        RECT 0.306 0.172 0.334 0.196 ;
        RECT 0.306 0.196 0.334 0.3827 ;
        RECT 0.306 0.3827 0.334 0.4013 ;
        RECT 0.334 0.0679 0.782 0.0867 ;
        RECT 0.782 0.0679 0.8139 0.0867 ;
        RECT 0.782 0.0867 0.8139 0.1533 ;
        RECT 0.782 0.1533 0.8139 0.1667 ;
        RECT 0.782 0.1667 0.8139 0.16678 ;
        RECT 0.782 0.172 0.8139 0.196 ;
        RECT 0.8139 0.1667 1.593 0.16678 ;
        RECT 0.8139 0.172 1.593 0.196 ;
  END
END TBUF_X12_8T

MACRO TBUF_X16_8T
  CLASS core ;
  FOREIGN TBUF_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.112 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.26 0.1419 0.324 ;
        RECT 0.114 0.324 0.1419 0.3427 ;
        RECT 0.1419 0.324 0.1739 0.3427 ;
        RECT 0.1739 0.324 0.24 0.3427 ;
        RECT 0.24 0.2133 0.272 0.26 ;
        RECT 0.24 0.26 0.272 0.324 ;
        RECT 0.24 0.324 0.272 0.3427 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.462 0.268 0.562 0.2987 ;
        RECT 0.562 0.2306 0.59 0.268 ;
        RECT 0.562 0.268 0.59 0.2987 ;
        RECT 0.59 0.268 0.6899 0.2987 ;
        RECT 0.6899 0.268 0.718 0.2987 ;
        RECT 0.6899 0.2987 0.718 0.384 ;
        RECT 0.718 0.268 0.902 0.2987 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.072 0.0427 1.104 0.0946 ;
        RECT 1.072 0.0946 1.104 0.1333 ;
        RECT 1.072 0.3467 1.104 0.384 ;
        RECT 1.072 0.384 1.104 0.4693 ;
        RECT 1.104 0.0946 1.968 0.1333 ;
        RECT 1.104 0.3467 1.968 0.384 ;
        RECT 1.968 0.0427 1.98 0.0946 ;
        RECT 1.968 0.0946 1.98 0.1333 ;
        RECT 1.968 0.3467 1.98 0.384 ;
        RECT 1.968 0.384 1.98 0.4693 ;
        RECT 1.98 0.0427 1.998 0.0946 ;
        RECT 1.98 0.0946 1.998 0.1333 ;
        RECT 1.98 0.3467 1.998 0.384 ;
        RECT 1.98 0.384 1.998 0.4693 ;
        RECT 1.998 0.0427 2 0.0946 ;
        RECT 1.998 0.0946 2 0.1333 ;
        RECT 1.998 0.3467 2 0.384 ;
        RECT 1.998 0.384 2 0.4693 ;
        RECT 2 0.0946 2.0339 0.1333 ;
        RECT 2 0.3467 2.0339 0.384 ;
        RECT 2.0339 0.0946 2.062 0.1333 ;
        RECT 2.0339 0.1333 2.062 0.3467 ;
        RECT 2.0339 0.3467 2.062 0.384 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.98 0.5307 ;
        RECT 1.98 0.4933 1.998 0.5307 ;
        RECT 1.998 0.4933 2.122 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 2.122 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.1747 ;
        RECT 0.05 0.1747 0.078 0.1933 ;
        RECT 0.05 0.1933 0.078 0.2306 ;
        RECT 0.05 0.2306 0.078 0.4 ;
        RECT 0.078 0.1747 0.1419 0.1933 ;
        RECT 0.1419 0.1747 0.1739 0.1933 ;
        RECT 0.1419 0.1933 0.1739 0.2306 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.398 0.132 ;
        RECT 0.274 0.4253 0.398 0.444 ;
        RECT 0.398 0.1107 0.426 0.132 ;
        RECT 0.398 0.132 0.426 0.2687 ;
        RECT 0.398 0.2687 0.426 0.3073 ;
        RECT 0.398 0.3073 0.426 0.4253 ;
        RECT 0.398 0.4253 0.426 0.444 ;
        RECT 0.426 0.4253 0.946 0.444 ;
        RECT 0.946 0.2687 0.974 0.3073 ;
        RECT 0.946 0.3073 0.974 0.4253 ;
        RECT 0.946 0.4253 0.974 0.444 ;
        RECT 0.974 0.2687 1.98 0.3073 ;
        RECT 0.146 0.3786 0.21 0.4013 ;
        RECT 0.21 0.0679 0.238 0.0867 ;
        RECT 0.21 0.0867 0.238 0.156 ;
        RECT 0.21 0.156 0.238 0.1747 ;
        RECT 0.21 0.3786 0.238 0.4013 ;
        RECT 0.238 0.0679 0.326 0.0867 ;
        RECT 0.238 0.156 0.326 0.1747 ;
        RECT 0.238 0.3786 0.326 0.4013 ;
        RECT 0.326 0.0679 0.362 0.0867 ;
        RECT 0.326 0.156 0.362 0.1747 ;
        RECT 0.326 0.1747 0.362 0.182 ;
        RECT 0.326 0.182 0.362 0.2207 ;
        RECT 0.326 0.2207 0.362 0.3786 ;
        RECT 0.326 0.3786 0.362 0.4013 ;
        RECT 0.362 0.0679 0.946 0.0867 ;
        RECT 0.946 0.0679 0.974 0.0867 ;
        RECT 0.946 0.0867 0.974 0.156 ;
        RECT 0.946 0.156 0.974 0.1747 ;
        RECT 0.946 0.1747 0.974 0.182 ;
        RECT 0.946 0.182 0.974 0.2207 ;
        RECT 0.974 0.182 1.998 0.2207 ;
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.1747 ;
        RECT 0.05 0.1747 0.078 0.1933 ;
        RECT 0.05 0.1933 0.078 0.2306 ;
        RECT 0.05 0.2306 0.078 0.4 ;
        RECT 0.078 0.1747 0.1419 0.1933 ;
        RECT 0.1419 0.1747 0.1739 0.1933 ;
        RECT 0.1419 0.1933 0.1739 0.2306 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.398 0.132 ;
        RECT 0.274 0.4253 0.398 0.444 ;
        RECT 0.398 0.1107 0.426 0.132 ;
        RECT 0.398 0.132 0.426 0.2687 ;
        RECT 0.398 0.2687 0.426 0.3073 ;
        RECT 0.398 0.3073 0.426 0.4253 ;
        RECT 0.398 0.4253 0.426 0.444 ;
        RECT 0.426 0.4253 0.946 0.444 ;
        RECT 0.946 0.2687 0.974 0.3073 ;
        RECT 0.946 0.3073 0.974 0.4253 ;
        RECT 0.946 0.4253 0.974 0.444 ;
        RECT 0.974 0.2687 1.98 0.3073 ;
        RECT 0.146 0.3786 0.21 0.4013 ;
        RECT 0.21 0.0679 0.238 0.0867 ;
        RECT 0.21 0.0867 0.238 0.156 ;
        RECT 0.21 0.156 0.238 0.1747 ;
        RECT 0.21 0.3786 0.238 0.4013 ;
        RECT 0.238 0.0679 0.326 0.0867 ;
        RECT 0.238 0.156 0.326 0.1747 ;
        RECT 0.238 0.3786 0.326 0.4013 ;
        RECT 0.326 0.0679 0.362 0.0867 ;
        RECT 0.326 0.156 0.362 0.1747 ;
        RECT 0.326 0.1747 0.362 0.182 ;
        RECT 0.326 0.182 0.362 0.2207 ;
        RECT 0.326 0.2207 0.362 0.3786 ;
        RECT 0.326 0.3786 0.362 0.4013 ;
        RECT 0.362 0.0679 0.946 0.0867 ;
        RECT 0.946 0.0679 0.974 0.0867 ;
        RECT 0.946 0.0867 0.974 0.156 ;
        RECT 0.946 0.156 0.974 0.1747 ;
        RECT 0.946 0.1747 0.974 0.182 ;
        RECT 0.946 0.182 0.974 0.2207 ;
        RECT 0.974 0.182 1.998 0.2207 ;
  END
END TBUF_X16_8T

MACRO TIEH_8T
  CLASS core ;
  FOREIGN TIEH_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.3153 0.1419 0.4693 ;
        RECT 0.1419 0.3153 0.147 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.202 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.202 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.064 0.1419 0.286 ;
      LAYER M1 ;
        RECT 0.114 0.064 0.1419 0.286 ;
  END
END TIEH_8T

MACRO TIEL_8T
  CLASS core ;
  FOREIGN TIEL_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.0427 0.147 0.1773 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.202 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.202 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.224 0.1419 0.448 ;
      LAYER M1 ;
        RECT 0.114 0.224 0.1419 0.448 ;
  END
END TIEL_8T

MACRO XNOR2_X1_8T
  CLASS core ;
  FOREIGN XNOR2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.168 0.21 0.1867 ;
        RECT 0.178 0.1867 0.21 0.2853 ;
        RECT 0.21 0.168 0.37 0.1867 ;
        RECT 0.37 0.168 0.398 0.1867 ;
        RECT 0.37 0.1867 0.398 0.2853 ;
        RECT 0.37 0.2853 0.398 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1613 0.078 0.2133 ;
        RECT 0.05 0.2133 0.078 0.4507 ;
        RECT 0.05 0.4507 0.078 0.4693 ;
        RECT 0.078 0.4507 0.274 0.4693 ;
        RECT 0.274 0.4507 0.498 0.4693 ;
        RECT 0.498 0.2133 0.526 0.4507 ;
        RECT 0.498 0.4507 0.526 0.4693 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.278 0.364 0.302 0.3647 ;
        RECT 0.278 0.3647 0.302 0.4007 ;
        RECT 0.278 0.4007 0.302 0.4013 ;
        RECT 0.302 0.1107 0.334 0.1293 ;
        RECT 0.302 0.364 0.334 0.3647 ;
        RECT 0.302 0.3647 0.334 0.4007 ;
        RECT 0.302 0.4007 0.334 0.4013 ;
        RECT 0.334 0.1107 0.434 0.1293 ;
        RECT 0.334 0.3647 0.434 0.4007 ;
        RECT 0.434 0.1107 0.462 0.1293 ;
        RECT 0.434 0.1653 0.462 0.184 ;
        RECT 0.434 0.184 0.462 0.364 ;
        RECT 0.434 0.364 0.462 0.3647 ;
        RECT 0.434 0.3647 0.462 0.4007 ;
        RECT 0.462 0.1107 0.493 0.1293 ;
        RECT 0.462 0.1653 0.493 0.184 ;
        RECT 0.493 0.1107 0.531 0.1293 ;
        RECT 0.493 0.1293 0.531 0.1653 ;
        RECT 0.493 0.1653 0.531 0.184 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.274 0.5307 ;
        RECT 0.274 0.4933 0.535 0.5307 ;
        RECT 0.535 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.0679 0.535 0.0867 ;
        RECT 0.114 0.1227 0.1419 0.144 ;
        RECT 0.114 0.144 0.1419 0.2267 ;
        RECT 0.114 0.2267 0.1419 0.3093 ;
        RECT 0.114 0.3093 0.1419 0.328 ;
        RECT 0.114 0.328 0.1419 0.368 ;
        RECT 0.1419 0.1227 0.234 0.144 ;
        RECT 0.1419 0.3093 0.234 0.328 ;
        RECT 0.234 0.3093 0.246 0.328 ;
        RECT 0.246 0.2267 0.274 0.3093 ;
        RECT 0.246 0.3093 0.274 0.328 ;
      LAYER M1 ;
        RECT 0.21 0.0679 0.535 0.0867 ;
        RECT 0.114 0.1227 0.1419 0.144 ;
        RECT 0.114 0.144 0.1419 0.2267 ;
        RECT 0.114 0.2267 0.1419 0.3093 ;
        RECT 0.114 0.3093 0.1419 0.328 ;
        RECT 0.114 0.328 0.1419 0.368 ;
        RECT 0.1419 0.1227 0.234 0.144 ;
        RECT 0.1419 0.3093 0.234 0.328 ;
        RECT 0.234 0.3093 0.246 0.328 ;
        RECT 0.246 0.2267 0.274 0.3093 ;
        RECT 0.246 0.3093 0.274 0.328 ;
  END
END XNOR2_X1_8T

MACRO XOR2_X1_8T
  CLASS core ;
  FOREIGN XOR2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.2293 0.21 0.324 ;
        RECT 0.178 0.324 0.21 0.3427 ;
        RECT 0.21 0.324 0.274 0.3427 ;
        RECT 0.274 0.324 0.37 0.3427 ;
        RECT 0.37 0.2133 0.398 0.2293 ;
        RECT 0.37 0.2293 0.398 0.324 ;
        RECT 0.37 0.324 0.398 0.3427 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0427 0.078 0.0613 ;
        RECT 0.05 0.0613 0.078 0.2987 ;
        RECT 0.05 0.2987 0.078 0.3507 ;
        RECT 0.078 0.0427 0.498 0.0613 ;
        RECT 0.498 0.0427 0.526 0.0613 ;
        RECT 0.498 0.0613 0.526 0.2987 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.275 0.1087 0.315 0.1093 ;
        RECT 0.275 0.1093 0.315 0.148 ;
        RECT 0.315 0.1087 0.334 0.1093 ;
        RECT 0.315 0.1093 0.334 0.148 ;
        RECT 0.315 0.3827 0.334 0.4013 ;
        RECT 0.334 0.1093 0.434 0.148 ;
        RECT 0.334 0.3827 0.434 0.4013 ;
        RECT 0.434 0.1093 0.462 0.148 ;
        RECT 0.434 0.148 0.462 0.328 ;
        RECT 0.434 0.328 0.462 0.3467 ;
        RECT 0.434 0.3827 0.462 0.4013 ;
        RECT 0.462 0.328 0.496 0.3467 ;
        RECT 0.462 0.3827 0.496 0.4013 ;
        RECT 0.496 0.328 0.34678 0.3467 ;
        RECT 0.496 0.3467 0.34678 0.3827 ;
        RECT 0.496 0.3827 0.528 0.4013 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.535 0.5307 ;
        RECT 0.535 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.246 0.4253 0.535 0.444 ;
        RECT 0.114 0.0907 0.1419 0.1867 ;
        RECT 0.114 0.1867 0.1419 0.2053 ;
        RECT 0.114 0.2053 0.1419 0.288 ;
        RECT 0.114 0.288 0.1419 0.368 ;
        RECT 0.114 0.368 0.1419 0.3893 ;
        RECT 0.1419 0.1867 0.246 0.2053 ;
        RECT 0.1419 0.368 0.246 0.3893 ;
        RECT 0.246 0.1867 0.247 0.2053 ;
        RECT 0.246 0.2053 0.247 0.288 ;
        RECT 0.246 0.368 0.247 0.3893 ;
        RECT 0.247 0.1867 0.274 0.2053 ;
        RECT 0.247 0.2053 0.274 0.288 ;
      LAYER M1 ;
        RECT 0.246 0.4253 0.535 0.444 ;
        RECT 0.114 0.0907 0.1419 0.1867 ;
        RECT 0.114 0.1867 0.1419 0.2053 ;
        RECT 0.114 0.2053 0.1419 0.288 ;
        RECT 0.114 0.288 0.1419 0.368 ;
        RECT 0.114 0.368 0.1419 0.3893 ;
        RECT 0.1419 0.1867 0.246 0.2053 ;
        RECT 0.1419 0.368 0.246 0.3893 ;
        RECT 0.246 0.1867 0.247 0.2053 ;
        RECT 0.246 0.2053 0.247 0.288 ;
        RECT 0.246 0.368 0.247 0.3893 ;
        RECT 0.247 0.1867 0.274 0.2053 ;
        RECT 0.247 0.2053 0.274 0.288 ;
  END
END XOR2_X1_8T

MACRO AND2_X1_12T
  CLASS core ;
  FOREIGN AND2_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.6959 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.127 0.078 0.525 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.114 0.334 0.64 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.162 0.1419 0.19 ;
        RECT 0.114 0.19 0.1419 0.428 ;
        RECT 0.114 0.428 0.1419 0.544 ;
        RECT 0.1419 0.162 0.242 0.19 ;
        RECT 0.242 0.162 0.27 0.19 ;
        RECT 0.242 0.19 0.27 0.428 ;
      LAYER M1 ;
        RECT 0.114 0.162 0.1419 0.19 ;
        RECT 0.114 0.19 0.1419 0.428 ;
        RECT 0.114 0.428 0.1419 0.544 ;
        RECT 0.1419 0.162 0.242 0.19 ;
        RECT 0.242 0.162 0.27 0.19 ;
        RECT 0.242 0.19 0.27 0.428 ;
  END
END AND2_X1_12T

MACRO AND2_X2_12T
  CLASS core ;
  FOREIGN AND2_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.672 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.248 0.083 0.52 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.064 0.306 0.13 ;
        RECT 0.302 0.638 0.306 0.704 ;
        RECT 0.306 0.064 0.334 0.13 ;
        RECT 0.306 0.13 0.334 0.638 ;
        RECT 0.306 0.638 0.334 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.574 0.082 0.602 ;
        RECT 0.082 0.166 0.242 0.194 ;
        RECT 0.082 0.574 0.242 0.602 ;
        RECT 0.242 0.166 0.27 0.194 ;
        RECT 0.242 0.194 0.27 0.574 ;
        RECT 0.242 0.574 0.27 0.602 ;
      LAYER M1 ;
        RECT 0.054 0.574 0.082 0.602 ;
        RECT 0.082 0.166 0.242 0.194 ;
        RECT 0.082 0.574 0.242 0.602 ;
        RECT 0.242 0.166 0.27 0.194 ;
        RECT 0.242 0.194 0.27 0.574 ;
        RECT 0.242 0.574 0.27 0.602 ;
  END
END AND2_X2_12T

MACRO AND3_X1_12T
  CLASS core ;
  FOREIGN AND3_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1729 0.192 0.211 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.192 0.08 0.576 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.114 0.462 0.654 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.079 0.1 0.238 0.132 ;
        RECT 0.054 0.631 0.274 0.659 ;
        RECT 0.274 0.095 0.37 0.137 ;
        RECT 0.274 0.631 0.37 0.659 ;
        RECT 0.37 0.095 0.398 0.137 ;
        RECT 0.37 0.137 0.398 0.631 ;
        RECT 0.37 0.631 0.398 0.659 ;
      LAYER M1 ;
        RECT 0.079 0.1 0.238 0.132 ;
        RECT 0.054 0.631 0.274 0.659 ;
        RECT 0.274 0.095 0.37 0.137 ;
        RECT 0.274 0.631 0.37 0.659 ;
        RECT 0.37 0.095 0.398 0.137 ;
        RECT 0.37 0.137 0.398 0.631 ;
        RECT 0.37 0.631 0.398 0.659 ;
  END
END AND3_X1_12T

MACRO AND3_X2_12T
  CLASS core ;
  FOREIGN AND3_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.32 0.206 0.513 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.256 0.083 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.302 0.27 0.537 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.366 0.064 0.37 0.157 ;
        RECT 0.366 0.638 0.37 0.704 ;
        RECT 0.37 0.064 0.398 0.157 ;
        RECT 0.37 0.157 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.072 0.08 0.156 ;
        RECT 0.048 0.156 0.08 0.188 ;
        RECT 0.08 0.156 0.298 0.188 ;
        RECT 0.054 0.581 0.146 0.613 ;
        RECT 0.146 0.224 0.306 0.252 ;
        RECT 0.146 0.581 0.306 0.613 ;
        RECT 0.306 0.224 0.334 0.252 ;
        RECT 0.306 0.252 0.334 0.581 ;
        RECT 0.306 0.581 0.334 0.613 ;
      LAYER M1 ;
        RECT 0.048 0.072 0.08 0.156 ;
        RECT 0.048 0.156 0.08 0.188 ;
        RECT 0.08 0.156 0.298 0.188 ;
        RECT 0.054 0.581 0.146 0.613 ;
        RECT 0.146 0.224 0.306 0.252 ;
        RECT 0.146 0.581 0.306 0.613 ;
        RECT 0.306 0.224 0.334 0.252 ;
        RECT 0.306 0.252 0.334 0.581 ;
        RECT 0.306 0.581 0.334 0.613 ;
  END
END AND3_X2_12T

MACRO AND4_X1_12T
  CLASS core ;
  FOREIGN AND4_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.192 0.272 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.1419 0.512 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.114 0.526 0.654 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.462 0.796 ;
        RECT 0.462 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.636 0.338 0.668 ;
        RECT 0.338 0.1 0.434 0.132 ;
        RECT 0.338 0.636 0.434 0.668 ;
        RECT 0.434 0.1 0.462 0.132 ;
        RECT 0.434 0.132 0.462 0.636 ;
        RECT 0.434 0.636 0.462 0.668 ;
        RECT 0.1409 0.099 0.298 0.147 ;
      LAYER M1 ;
        RECT 0.082 0.636 0.338 0.668 ;
        RECT 0.338 0.1 0.434 0.132 ;
        RECT 0.338 0.636 0.434 0.668 ;
        RECT 0.434 0.1 0.462 0.132 ;
        RECT 0.434 0.132 0.462 0.636 ;
        RECT 0.434 0.636 0.462 0.668 ;
        RECT 0.1409 0.099 0.298 0.147 ;
  END
END AND4_X1_12T

MACRO AND4_X2_12T
  CLASS core ;
  FOREIGN AND4_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.96 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.241 0.398 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.192 0.27 0.577 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.1419 0.577 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.577 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.096 0.526 0.64 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.462 0.796 ;
        RECT 0.462 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.1419 0.1 0.298 0.132 ;
        RECT 0.082 0.636 0.342 0.668 ;
        RECT 0.342 0.165 0.434 0.197 ;
        RECT 0.342 0.636 0.434 0.668 ;
        RECT 0.434 0.165 0.462 0.197 ;
        RECT 0.434 0.197 0.462 0.636 ;
        RECT 0.434 0.636 0.462 0.668 ;
      LAYER M1 ;
        RECT 0.1419 0.1 0.298 0.132 ;
        RECT 0.082 0.636 0.342 0.668 ;
        RECT 0.342 0.165 0.434 0.197 ;
        RECT 0.342 0.636 0.434 0.668 ;
        RECT 0.434 0.165 0.462 0.197 ;
        RECT 0.434 0.197 0.462 0.636 ;
        RECT 0.434 0.636 0.462 0.668 ;
  END
END AND4_X2_12T

MACRO ANTENNA_12T
  CLASS core ;
  FOREIGN ANTENNA_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.288 BY 0.512 ;
END ANTENNA_12T

MACRO AOI21_X1_12T
  CLASS core ;
  FOREIGN AOI21_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.192 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.134 0.078 0.512 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.512 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1 0.1419 0.132 ;
        RECT 0.114 0.132 0.1419 0.536 ;
        RECT 0.1419 0.1 0.306 0.132 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.298 0.796 ;
        RECT 0.298 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.58 0.08 0.612 ;
        RECT 0.048 0.612 0.08 0.704 ;
        RECT 0.08 0.58 0.298 0.612 ;
      LAYER M1 ;
        RECT 0.048 0.58 0.08 0.612 ;
        RECT 0.048 0.612 0.08 0.704 ;
        RECT 0.08 0.58 0.298 0.612 ;
  END
END AOI21_X1_12T

MACRO AOI21_X2_12T
  CLASS core ;
  FOREIGN AOI21_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.302 0.398 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.23 0.27 0.258 ;
        RECT 0.242 0.258 0.27 0.448 ;
        RECT 0.242 0.448 0.27 0.512 ;
        RECT 0.27 0.23 0.493 0.258 ;
        RECT 0.493 0.23 0.531 0.258 ;
        RECT 0.493 0.258 0.531 0.448 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.448 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.077 0.166 0.178 0.194 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.489 ;
        RECT 0.178 0.489 0.206 0.5709 ;
        RECT 0.178 0.5709 0.206 0.599 ;
        RECT 0.206 0.166 0.43 0.194 ;
        RECT 0.206 0.5709 0.43 0.599 ;
        RECT 0.43 0.5709 0.434 0.599 ;
        RECT 0.434 0.489 0.462 0.5709 ;
        RECT 0.434 0.5709 0.462 0.599 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.535 0.796 ;
        RECT 0.535 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.55 0.08 0.635 ;
        RECT 0.048 0.635 0.08 0.669 ;
        RECT 0.08 0.635 0.498 0.669 ;
        RECT 0.498 0.516 0.526 0.55 ;
        RECT 0.498 0.55 0.526 0.635 ;
        RECT 0.498 0.635 0.526 0.669 ;
        RECT 0.146 0.1019 0.535 0.13 ;
      LAYER M1 ;
        RECT 0.048 0.55 0.08 0.635 ;
        RECT 0.048 0.635 0.08 0.669 ;
        RECT 0.08 0.635 0.498 0.669 ;
        RECT 0.498 0.516 0.526 0.55 ;
        RECT 0.498 0.55 0.526 0.635 ;
        RECT 0.498 0.635 0.526 0.669 ;
        RECT 0.146 0.1019 0.535 0.13 ;
  END
END AOI21_X2_12T

MACRO AOI22_X1_12T
  CLASS core ;
  FOREIGN AOI22_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.672 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.192 0.27 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.485 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.198 0.1419 0.576 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1409 0.1019 0.306 0.13 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.13 0.334 0.582 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.63 0.37 0.674 ;
        RECT 0.37 0.553 0.398 0.63 ;
        RECT 0.37 0.63 0.398 0.674 ;
      LAYER M1 ;
        RECT 0.082 0.63 0.37 0.674 ;
        RECT 0.37 0.553 0.398 0.63 ;
        RECT 0.37 0.63 0.398 0.674 ;
  END
END AOI22_X1_12T

MACRO AOI22_X2_12T
  CLASS core ;
  FOREIGN AOI22_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.152 BY 1.152 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.274 0.462 0.302 ;
        RECT 0.434 0.302 0.462 0.489 ;
        RECT 0.434 0.489 0.462 0.512 ;
        RECT 0.462 0.274 0.654 0.302 ;
        RECT 0.654 0.274 0.6899 0.302 ;
        RECT 0.6899 0.274 0.718 0.302 ;
        RECT 0.6899 0.302 0.718 0.489 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.37 0.59 0.512 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.306 0.334 0.526 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.242 0.078 0.512 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2 0.27 0.228 ;
        RECT 0.242 0.228 0.27 0.229 ;
        RECT 0.242 0.229 0.27 0.32 ;
        RECT 0.27 0.2 0.362 0.228 ;
        RECT 0.362 0.2 0.37 0.228 ;
        RECT 0.37 0.2 0.398 0.228 ;
        RECT 0.37 0.228 0.398 0.229 ;
        RECT 0.37 0.229 0.398 0.32 ;
        RECT 0.37 0.32 0.398 0.463 ;
        RECT 0.37 0.463 0.398 0.5679 ;
        RECT 0.37 0.5679 0.398 0.602 ;
        RECT 0.398 0.2 0.626 0.228 ;
        RECT 0.398 0.228 0.626 0.229 ;
        RECT 0.398 0.5679 0.626 0.602 ;
        RECT 0.626 0.2 0.654 0.228 ;
        RECT 0.626 0.228 0.654 0.229 ;
        RECT 0.626 0.463 0.654 0.5679 ;
        RECT 0.626 0.5679 0.654 0.602 ;
        RECT 0.654 0.2 0.6899 0.228 ;
        RECT 0.654 0.228 0.6899 0.229 ;
        RECT 0.6899 0.096 0.718 0.2 ;
        RECT 0.6899 0.2 0.718 0.228 ;
        RECT 0.6899 0.228 0.718 0.229 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.718 0.796 ;
        RECT 0.718 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.406 0.132 0.626 0.164 ;
        RECT 0.626 0.072 0.654 0.132 ;
        RECT 0.626 0.132 0.654 0.164 ;
        RECT 0.077 0.638 0.6899 0.666 ;
        RECT 0.6899 0.557 0.718 0.638 ;
        RECT 0.6899 0.638 0.718 0.666 ;
        RECT 0.0859 0.0869 0.362 0.145 ;
      LAYER M1 ;
        RECT 0.406 0.132 0.626 0.164 ;
        RECT 0.626 0.072 0.654 0.132 ;
        RECT 0.626 0.132 0.654 0.164 ;
        RECT 0.077 0.638 0.6899 0.666 ;
        RECT 0.6899 0.557 0.718 0.638 ;
        RECT 0.6899 0.638 0.718 0.666 ;
        RECT 0.0859 0.0869 0.362 0.145 ;
  END
END AOI22_X2_12T

MACRO BUF_X1_12T
  CLASS core ;
  FOREIGN BUF_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.48 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.114 0.272 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1429 0.796 ;
        RECT 0.1429 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.072 0.115 0.185 ;
        RECT 0.114 0.185 0.115 0.213 ;
        RECT 0.114 0.428 0.115 0.456 ;
        RECT 0.114 0.456 0.115 0.558 ;
        RECT 0.115 0.072 0.1419 0.185 ;
        RECT 0.115 0.185 0.1419 0.213 ;
        RECT 0.115 0.213 0.1419 0.428 ;
        RECT 0.115 0.428 0.1419 0.456 ;
        RECT 0.115 0.456 0.1419 0.558 ;
        RECT 0.1419 0.185 0.1429 0.213 ;
        RECT 0.1419 0.213 0.1429 0.428 ;
        RECT 0.1419 0.428 0.1429 0.456 ;
      LAYER M1 ;
        RECT 0.114 0.072 0.115 0.185 ;
        RECT 0.114 0.185 0.115 0.213 ;
        RECT 0.114 0.428 0.115 0.456 ;
        RECT 0.114 0.456 0.115 0.558 ;
        RECT 0.115 0.072 0.1419 0.185 ;
        RECT 0.115 0.185 0.1419 0.213 ;
        RECT 0.115 0.213 0.1419 0.428 ;
        RECT 0.115 0.428 0.1419 0.456 ;
        RECT 0.115 0.456 0.1419 0.558 ;
        RECT 0.1419 0.185 0.1429 0.213 ;
        RECT 0.1419 0.213 0.1429 0.428 ;
        RECT 0.1419 0.428 0.1429 0.456 ;
  END
END BUF_X1_12T

MACRO BUF_X2_12T
  CLASS core ;
  FOREIGN BUF_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.48 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.267 0.078 0.512 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1739 0.603 0.177 0.704 ;
        RECT 0.177 0.072 0.178 0.132 ;
        RECT 0.177 0.603 0.178 0.704 ;
        RECT 0.178 0.072 0.206 0.132 ;
        RECT 0.178 0.132 0.206 0.603 ;
        RECT 0.178 0.603 0.206 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.042 0.556 0.05 0.584 ;
        RECT 0.042 0.584 0.05 0.686 ;
        RECT 0.05 0.096 0.078 0.192 ;
        RECT 0.05 0.192 0.078 0.22 ;
        RECT 0.05 0.556 0.078 0.584 ;
        RECT 0.05 0.584 0.078 0.686 ;
        RECT 0.078 0.192 0.0859 0.22 ;
        RECT 0.078 0.556 0.0859 0.584 ;
        RECT 0.078 0.584 0.0859 0.686 ;
        RECT 0.0859 0.192 0.114 0.22 ;
        RECT 0.0859 0.556 0.114 0.584 ;
        RECT 0.114 0.192 0.1419 0.22 ;
        RECT 0.114 0.22 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
      LAYER M1 ;
        RECT 0.042 0.556 0.05 0.584 ;
        RECT 0.042 0.584 0.05 0.686 ;
        RECT 0.05 0.096 0.078 0.192 ;
        RECT 0.05 0.192 0.078 0.22 ;
        RECT 0.05 0.556 0.078 0.584 ;
        RECT 0.05 0.584 0.078 0.686 ;
        RECT 0.078 0.192 0.0859 0.22 ;
        RECT 0.078 0.556 0.0859 0.584 ;
        RECT 0.078 0.584 0.0859 0.686 ;
        RECT 0.0859 0.192 0.114 0.22 ;
        RECT 0.0859 0.556 0.114 0.584 ;
        RECT 0.114 0.192 0.1419 0.22 ;
        RECT 0.114 0.22 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
  END
END BUF_X2_12T

MACRO BUF_X4_12T
  CLASS core ;
  FOREIGN BUF_X4_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.242 0.206 0.526 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.1019 0.21 0.13 ;
        RECT 0.21 0.1019 0.27 0.13 ;
        RECT 0.21 0.638 0.27 0.666 ;
        RECT 0.27 0.1019 0.368 0.13 ;
        RECT 0.27 0.638 0.368 0.666 ;
        RECT 0.368 0.1019 0.4 0.13 ;
        RECT 0.368 0.13 0.4 0.638 ;
        RECT 0.368 0.638 0.4 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.027 0.166 0.0859 0.198 ;
        RECT 0.0859 0.166 0.242 0.198 ;
        RECT 0.0859 0.5699 0.242 0.602 ;
        RECT 0.242 0.166 0.27 0.198 ;
        RECT 0.242 0.198 0.27 0.5699 ;
        RECT 0.242 0.5699 0.27 0.602 ;
      LAYER M1 ;
        RECT 0.027 0.166 0.0859 0.198 ;
        RECT 0.0859 0.166 0.242 0.198 ;
        RECT 0.0859 0.5699 0.242 0.602 ;
        RECT 0.242 0.166 0.27 0.198 ;
        RECT 0.242 0.198 0.27 0.5699 ;
        RECT 0.242 0.5699 0.27 0.602 ;
  END
END BUF_X4_12T

MACRO BUF_X8_12T
  CLASS core ;
  FOREIGN BUF_X8_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.344 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.366 ;
        RECT 0.05 0.366 0.078 0.398 ;
        RECT 0.05 0.398 0.078 0.512 ;
        RECT 0.078 0.366 0.298 0.398 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.1019 0.7 0.13 ;
        RECT 0.338 0.638 0.7 0.666 ;
        RECT 0.7 0.1019 0.754 0.13 ;
        RECT 0.7 0.638 0.754 0.666 ;
        RECT 0.754 0.1019 0.782 0.13 ;
        RECT 0.754 0.13 0.782 0.638 ;
        RECT 0.754 0.638 0.782 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.7 0.796 ;
        RECT 0.7 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.099 0.098 0.114 0.186 ;
        RECT 0.099 0.186 0.114 0.214 ;
        RECT 0.114 0.098 0.1419 0.186 ;
        RECT 0.114 0.186 0.1419 0.214 ;
        RECT 0.114 0.527 0.1419 0.583 ;
        RECT 0.114 0.583 0.1419 0.67 ;
        RECT 0.1419 0.098 0.157 0.186 ;
        RECT 0.1419 0.186 0.157 0.214 ;
        RECT 0.1419 0.527 0.157 0.583 ;
        RECT 0.157 0.186 0.354 0.214 ;
        RECT 0.157 0.527 0.354 0.583 ;
        RECT 0.354 0.186 0.382 0.214 ;
        RECT 0.354 0.214 0.382 0.341 ;
        RECT 0.354 0.341 0.382 0.369 ;
        RECT 0.354 0.369 0.382 0.527 ;
        RECT 0.354 0.527 0.382 0.583 ;
        RECT 0.382 0.341 0.7 0.369 ;
      LAYER M1 ;
        RECT 0.099 0.098 0.114 0.186 ;
        RECT 0.099 0.186 0.114 0.214 ;
        RECT 0.114 0.098 0.1419 0.186 ;
        RECT 0.114 0.186 0.1419 0.214 ;
        RECT 0.114 0.527 0.1419 0.583 ;
        RECT 0.114 0.583 0.1419 0.67 ;
        RECT 0.1419 0.098 0.157 0.186 ;
        RECT 0.1419 0.186 0.157 0.214 ;
        RECT 0.1419 0.527 0.157 0.583 ;
        RECT 0.157 0.186 0.354 0.214 ;
        RECT 0.157 0.527 0.354 0.583 ;
        RECT 0.354 0.186 0.382 0.214 ;
        RECT 0.354 0.214 0.382 0.341 ;
        RECT 0.354 0.341 0.382 0.369 ;
        RECT 0.354 0.369 0.382 0.527 ;
        RECT 0.354 0.527 0.382 0.583 ;
        RECT 0.382 0.341 0.7 0.369 ;
  END
END BUF_X8_12T

MACRO BUF_X12_12T
  CLASS core ;
  FOREIGN BUF_X12_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.92 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.236 0.08 0.366 ;
        RECT 0.048 0.366 0.08 0.398 ;
        RECT 0.048 0.398 0.08 0.515 ;
        RECT 0.08 0.366 0.426 0.398 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.1019 1.07 0.13 ;
        RECT 0.466 0.638 1.07 0.666 ;
        RECT 1.07 0.1019 1.1359 0.13 ;
        RECT 1.07 0.638 1.1359 0.666 ;
        RECT 1.1359 0.1019 1.168 0.13 ;
        RECT 1.1359 0.13 1.168 0.638 ;
        RECT 1.1359 0.638 1.168 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.07 0.796 ;
        RECT 1.07 0.74 1.29 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.29 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.098 0.551 0.112 0.583 ;
        RECT 0.098 0.583 0.112 0.67 ;
        RECT 0.112 0.098 0.144 0.185 ;
        RECT 0.112 0.185 0.144 0.217 ;
        RECT 0.112 0.551 0.144 0.583 ;
        RECT 0.112 0.583 0.144 0.67 ;
        RECT 0.144 0.185 0.157 0.217 ;
        RECT 0.144 0.551 0.157 0.583 ;
        RECT 0.144 0.583 0.157 0.67 ;
        RECT 0.157 0.185 0.462 0.217 ;
        RECT 0.157 0.551 0.462 0.583 ;
        RECT 0.462 0.185 0.49 0.217 ;
        RECT 0.462 0.217 0.49 0.37 ;
        RECT 0.462 0.37 0.49 0.398 ;
        RECT 0.462 0.398 0.49 0.551 ;
        RECT 0.462 0.551 0.49 0.583 ;
        RECT 0.49 0.37 1.07 0.398 ;
      LAYER M1 ;
        RECT 0.098 0.551 0.112 0.583 ;
        RECT 0.098 0.583 0.112 0.67 ;
        RECT 0.112 0.098 0.144 0.185 ;
        RECT 0.112 0.185 0.144 0.217 ;
        RECT 0.112 0.551 0.144 0.583 ;
        RECT 0.112 0.583 0.144 0.67 ;
        RECT 0.144 0.185 0.157 0.217 ;
        RECT 0.144 0.551 0.157 0.583 ;
        RECT 0.144 0.583 0.157 0.67 ;
        RECT 0.157 0.185 0.462 0.217 ;
        RECT 0.157 0.551 0.462 0.583 ;
        RECT 0.462 0.185 0.49 0.217 ;
        RECT 0.462 0.217 0.49 0.37 ;
        RECT 0.462 0.37 0.49 0.398 ;
        RECT 0.462 0.398 0.49 0.551 ;
        RECT 0.462 0.551 0.49 0.583 ;
        RECT 0.49 0.37 1.07 0.398 ;
  END
END BUF_X12_12T

MACRO BUF_X16_12T
  CLASS core ;
  FOREIGN BUF_X16_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.496 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.232 0.078 0.355 ;
        RECT 0.05 0.355 0.078 0.413 ;
        RECT 0.05 0.413 0.078 0.512 ;
        RECT 0.078 0.355 0.554 0.413 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.1019 1.454 0.13 ;
        RECT 0.594 0.632 1.454 0.66 ;
        RECT 1.454 0.1019 1.52 0.13 ;
        RECT 1.454 0.632 1.52 0.66 ;
        RECT 1.52 0.1019 1.552 0.13 ;
        RECT 1.52 0.13 1.552 0.632 ;
        RECT 1.52 0.632 1.552 0.66 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.454 0.796 ;
        RECT 1.454 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.098 0.1419 0.205 ;
        RECT 0.114 0.205 0.1419 0.233 ;
        RECT 0.114 0.458 0.1419 0.486 ;
        RECT 0.114 0.486 0.1419 0.643 ;
        RECT 0.1419 0.205 0.59 0.233 ;
        RECT 0.1419 0.458 0.59 0.486 ;
        RECT 0.59 0.205 0.618 0.233 ;
        RECT 0.59 0.233 0.618 0.368 ;
        RECT 0.59 0.368 0.618 0.396 ;
        RECT 0.59 0.396 0.618 0.458 ;
        RECT 0.59 0.458 0.618 0.486 ;
        RECT 0.618 0.368 1.454 0.396 ;
      LAYER M1 ;
        RECT 0.114 0.098 0.1419 0.205 ;
        RECT 0.114 0.205 0.1419 0.233 ;
        RECT 0.114 0.458 0.1419 0.486 ;
        RECT 0.114 0.486 0.1419 0.643 ;
        RECT 0.1419 0.205 0.59 0.233 ;
        RECT 0.1419 0.458 0.59 0.486 ;
        RECT 0.59 0.205 0.618 0.233 ;
        RECT 0.59 0.233 0.618 0.368 ;
        RECT 0.59 0.368 0.618 0.396 ;
        RECT 0.59 0.396 0.618 0.458 ;
        RECT 0.59 0.458 0.618 0.486 ;
        RECT 0.618 0.368 1.454 0.396 ;
  END
END BUF_X16_12T

MACRO CLKBUF_X1_12T
  CLASS core ;
  FOREIGN CLKBUF_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.48 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.114 0.272 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1429 0.796 ;
        RECT 0.1429 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.072 0.115 0.185 ;
        RECT 0.114 0.185 0.115 0.213 ;
        RECT 0.114 0.393 0.115 0.458 ;
        RECT 0.114 0.458 0.115 0.523 ;
        RECT 0.115 0.072 0.1419 0.185 ;
        RECT 0.115 0.185 0.1419 0.213 ;
        RECT 0.115 0.213 0.1419 0.393 ;
        RECT 0.115 0.393 0.1419 0.458 ;
        RECT 0.115 0.458 0.1419 0.523 ;
        RECT 0.1419 0.185 0.1429 0.213 ;
        RECT 0.1419 0.213 0.1429 0.393 ;
        RECT 0.1419 0.393 0.1429 0.458 ;
      LAYER M1 ;
        RECT 0.114 0.072 0.115 0.185 ;
        RECT 0.114 0.185 0.115 0.213 ;
        RECT 0.114 0.393 0.115 0.458 ;
        RECT 0.114 0.458 0.115 0.523 ;
        RECT 0.115 0.072 0.1419 0.185 ;
        RECT 0.115 0.185 0.1419 0.213 ;
        RECT 0.115 0.213 0.1419 0.393 ;
        RECT 0.115 0.393 0.1419 0.458 ;
        RECT 0.115 0.458 0.1419 0.523 ;
        RECT 0.1419 0.185 0.1429 0.213 ;
        RECT 0.1419 0.213 0.1429 0.393 ;
        RECT 0.1419 0.393 0.1429 0.458 ;
  END
END CLKBUF_X1_12T

MACRO CLKBUF_X2_12T
  CLASS core ;
  FOREIGN CLKBUF_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.48 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.296 0.078 0.512 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1739 0.638 0.178 0.704 ;
        RECT 0.178 0.072 0.206 0.638 ;
        RECT 0.178 0.638 0.206 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.129 0.08 0.192 ;
        RECT 0.048 0.192 0.08 0.22 ;
        RECT 0.048 0.556 0.08 0.584 ;
        RECT 0.048 0.584 0.08 0.686 ;
        RECT 0.08 0.192 0.114 0.22 ;
        RECT 0.08 0.556 0.114 0.584 ;
        RECT 0.114 0.192 0.1419 0.22 ;
        RECT 0.114 0.22 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
      LAYER M1 ;
        RECT 0.048 0.129 0.08 0.192 ;
        RECT 0.048 0.192 0.08 0.22 ;
        RECT 0.048 0.556 0.08 0.584 ;
        RECT 0.048 0.584 0.08 0.686 ;
        RECT 0.08 0.192 0.114 0.22 ;
        RECT 0.08 0.556 0.114 0.584 ;
        RECT 0.114 0.192 0.1419 0.22 ;
        RECT 0.114 0.22 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
  END
END CLKBUF_X2_12T

MACRO CLKBUF_X4_12T
  CLASS core ;
  FOREIGN CLKBUF_X4_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.1419 0.526 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.1019 0.205 0.13 ;
        RECT 0.205 0.1019 0.206 0.13 ;
        RECT 0.205 0.638 0.206 0.666 ;
        RECT 0.206 0.1019 0.368 0.13 ;
        RECT 0.206 0.638 0.368 0.666 ;
        RECT 0.368 0.1019 0.4 0.13 ;
        RECT 0.368 0.13 0.4 0.638 ;
        RECT 0.368 0.638 0.4 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.041 0.166 0.082 0.194 ;
        RECT 0.082 0.166 0.178 0.194 ;
        RECT 0.082 0.574 0.178 0.602 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.574 ;
        RECT 0.178 0.574 0.206 0.602 ;
      LAYER M1 ;
        RECT 0.041 0.166 0.082 0.194 ;
        RECT 0.082 0.166 0.178 0.194 ;
        RECT 0.082 0.574 0.178 0.602 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.574 ;
        RECT 0.178 0.574 0.206 0.602 ;
  END
END CLKBUF_X4_12T

MACRO CLKBUF_X8_12T
  CLASS core ;
  FOREIGN CLKBUF_X8_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.344 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.328 ;
        RECT 0.05 0.328 0.078 0.356 ;
        RECT 0.05 0.356 0.078 0.512 ;
        RECT 0.078 0.256 0.079 0.328 ;
        RECT 0.078 0.328 0.079 0.356 ;
        RECT 0.079 0.328 0.318 0.356 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.1019 0.718 0.13 ;
        RECT 0.338 0.638 0.718 0.666 ;
        RECT 0.718 0.1019 0.754 0.13 ;
        RECT 0.718 0.638 0.754 0.666 ;
        RECT 0.754 0.1019 0.782 0.13 ;
        RECT 0.754 0.13 0.782 0.638 ;
        RECT 0.754 0.638 0.782 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.718 0.796 ;
        RECT 0.718 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.166 0.114 0.194 ;
        RECT 0.114 0.166 0.1419 0.194 ;
        RECT 0.114 0.45 0.1419 0.482 ;
        RECT 0.114 0.482 0.1419 0.542 ;
        RECT 0.1419 0.166 0.406 0.194 ;
        RECT 0.1419 0.45 0.406 0.482 ;
        RECT 0.406 0.166 0.434 0.194 ;
        RECT 0.406 0.194 0.434 0.357 ;
        RECT 0.406 0.357 0.434 0.415 ;
        RECT 0.406 0.415 0.434 0.45 ;
        RECT 0.406 0.45 0.434 0.482 ;
        RECT 0.434 0.357 0.718 0.415 ;
      LAYER M1 ;
        RECT 0.05 0.166 0.114 0.194 ;
        RECT 0.114 0.166 0.1419 0.194 ;
        RECT 0.114 0.45 0.1419 0.482 ;
        RECT 0.114 0.482 0.1419 0.542 ;
        RECT 0.1419 0.166 0.406 0.194 ;
        RECT 0.1419 0.45 0.406 0.482 ;
        RECT 0.406 0.166 0.434 0.194 ;
        RECT 0.406 0.194 0.434 0.357 ;
        RECT 0.406 0.357 0.434 0.415 ;
        RECT 0.406 0.415 0.434 0.45 ;
        RECT 0.406 0.45 0.434 0.482 ;
        RECT 0.434 0.357 0.718 0.415 ;
  END
END CLKBUF_X8_12T

MACRO CLKBUF_X12_12T
  CLASS core ;
  FOREIGN CLKBUF_X12_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.92 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.238 0.083 0.336 ;
        RECT 0.045 0.336 0.083 0.368 ;
        RECT 0.045 0.368 0.083 0.53 ;
        RECT 0.083 0.336 0.426 0.368 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.1019 0.998 0.13 ;
        RECT 0.466 0.638 0.998 0.666 ;
        RECT 0.998 0.1019 1.1359 0.13 ;
        RECT 0.998 0.638 1.1359 0.666 ;
        RECT 1.1359 0.1019 1.168 0.13 ;
        RECT 1.1359 0.13 1.168 0.638 ;
        RECT 1.1359 0.638 1.168 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.998 0.796 ;
        RECT 0.998 0.74 1.29 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.29 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0429 0.166 0.114 0.194 ;
        RECT 0.114 0.166 0.1419 0.194 ;
        RECT 0.114 0.55 0.1419 0.578 ;
        RECT 0.114 0.578 0.1419 0.67 ;
        RECT 0.1419 0.166 0.462 0.194 ;
        RECT 0.1419 0.55 0.462 0.578 ;
        RECT 0.462 0.166 0.49 0.194 ;
        RECT 0.462 0.194 0.49 0.314 ;
        RECT 0.462 0.314 0.49 0.3459 ;
        RECT 0.462 0.3459 0.49 0.55 ;
        RECT 0.462 0.55 0.49 0.578 ;
        RECT 0.49 0.166 0.494 0.194 ;
        RECT 0.49 0.194 0.494 0.314 ;
        RECT 0.49 0.314 0.494 0.3459 ;
        RECT 0.494 0.314 0.998 0.3459 ;
      LAYER M1 ;
        RECT 0.0429 0.166 0.114 0.194 ;
        RECT 0.114 0.166 0.1419 0.194 ;
        RECT 0.114 0.55 0.1419 0.578 ;
        RECT 0.114 0.578 0.1419 0.67 ;
        RECT 0.1419 0.166 0.462 0.194 ;
        RECT 0.1419 0.55 0.462 0.578 ;
        RECT 0.462 0.166 0.49 0.194 ;
        RECT 0.462 0.194 0.49 0.314 ;
        RECT 0.462 0.314 0.49 0.3459 ;
        RECT 0.462 0.3459 0.49 0.55 ;
        RECT 0.462 0.55 0.49 0.578 ;
        RECT 0.49 0.166 0.494 0.194 ;
        RECT 0.49 0.194 0.494 0.314 ;
        RECT 0.49 0.314 0.494 0.3459 ;
        RECT 0.494 0.314 0.998 0.3459 ;
  END
END CLKBUF_X12_12T

MACRO CLKBUF_X16_12T
  CLASS core ;
  FOREIGN CLKBUF_X16_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.496 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.222 0.078 0.326 ;
        RECT 0.05 0.326 0.078 0.358 ;
        RECT 0.05 0.358 0.078 0.526 ;
        RECT 0.078 0.326 0.554 0.358 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.0869 1.454 0.145 ;
        RECT 0.594 0.623 1.454 0.681 ;
        RECT 1.454 0.0869 1.52 0.145 ;
        RECT 1.454 0.623 1.52 0.681 ;
        RECT 1.52 0.0869 1.552 0.145 ;
        RECT 1.52 0.145 1.552 0.623 ;
        RECT 1.52 0.623 1.552 0.681 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.454 0.796 ;
        RECT 1.454 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.109 0.1419 0.205 ;
        RECT 0.114 0.205 0.1419 0.233 ;
        RECT 0.114 0.525 0.1419 0.5629 ;
        RECT 0.114 0.5629 0.1419 0.638 ;
        RECT 0.1419 0.205 0.595 0.233 ;
        RECT 0.1419 0.525 0.595 0.5629 ;
        RECT 0.595 0.205 0.653 0.233 ;
        RECT 0.595 0.233 0.653 0.316 ;
        RECT 0.595 0.316 0.653 0.3439 ;
        RECT 0.595 0.3439 0.653 0.525 ;
        RECT 0.595 0.525 0.653 0.5629 ;
        RECT 0.653 0.316 1.454 0.3439 ;
      LAYER M1 ;
        RECT 0.114 0.109 0.1419 0.205 ;
        RECT 0.114 0.205 0.1419 0.233 ;
        RECT 0.114 0.525 0.1419 0.5629 ;
        RECT 0.114 0.5629 0.1419 0.638 ;
        RECT 0.1419 0.205 0.595 0.233 ;
        RECT 0.1419 0.525 0.595 0.5629 ;
        RECT 0.595 0.205 0.653 0.233 ;
        RECT 0.595 0.233 0.653 0.316 ;
        RECT 0.595 0.316 0.653 0.3439 ;
        RECT 0.595 0.3439 0.653 0.525 ;
        RECT 0.595 0.525 0.653 0.5629 ;
        RECT 0.653 0.316 1.454 0.3439 ;
  END
END CLKBUF_X16_12T

MACRO CLKGATETST_X1_12T
  CLASS core ;
  FOREIGN CLKGATETST_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.632 BY 0.512 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.6899 0.238 0.718 0.512 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.672 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.32 0.078 0.672 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.01 0.096 1.038 0.654 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.366 0.796 ;
        RECT 0.366 0.74 0.91 0.796 ;
        RECT 0.91 0.74 0.974 0.796 ;
        RECT 0.974 0.74 1.098 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.098 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.21 0.402 0.686 0.43 ;
        RECT 0.146 0.466 0.522 0.494 ;
        RECT 0.73 0.402 1.006 0.43 ;
      LAYER MINT1 ;
        RECT 0.21 0.402 0.686 0.43 ;
        RECT 0.146 0.466 0.522 0.494 ;
        RECT 0.73 0.402 1.006 0.43 ;
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.238 0.13 ;
        RECT 0.242 0.264 0.27 0.541 ;
        RECT 0.37 0.242 0.398 0.502 ;
        RECT 0.462 0.372 0.494 0.51 ;
        RECT 0.626 0.166 0.654 0.194 ;
        RECT 0.626 0.194 0.654 0.556 ;
        RECT 0.626 0.556 0.654 0.592 ;
        RECT 0.654 0.166 0.75 0.194 ;
        RECT 0.654 0.556 0.75 0.592 ;
        RECT 0.75 0.166 0.755 0.194 ;
        RECT 0.754 0.248 0.79 0.463 ;
        RECT 0.754 0.463 0.79 0.502 ;
        RECT 0.79 0.463 0.8179 0.502 ;
        RECT 0.8179 0.463 0.846 0.502 ;
        RECT 0.8179 0.502 0.846 0.584 ;
        RECT 0.946 0.226 0.974 0.574 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.628 ;
        RECT 0.178 0.628 0.206 0.676 ;
        RECT 0.206 0.166 0.302 0.194 ;
        RECT 0.206 0.628 0.302 0.676 ;
        RECT 0.302 0.628 0.366 0.676 ;
        RECT 0.306 0.307 0.334 0.546 ;
        RECT 0.306 0.546 0.334 0.574 ;
        RECT 0.334 0.546 0.558 0.574 ;
        RECT 0.558 0.184 0.59 0.307 ;
        RECT 0.558 0.307 0.59 0.546 ;
        RECT 0.558 0.546 0.59 0.574 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.334 ;
        RECT 0.462 0.1019 0.466 0.13 ;
        RECT 0.466 0.1019 0.882 0.13 ;
        RECT 0.466 0.628 0.882 0.676 ;
        RECT 0.882 0.1019 0.91 0.13 ;
        RECT 0.882 0.13 0.91 0.334 ;
        RECT 0.882 0.334 0.91 0.628 ;
        RECT 0.882 0.628 0.91 0.676 ;
      LAYER V1 ;
        RECT 0.178 0.466 0.206 0.494 ;
        RECT 0.242 0.402 0.27 0.43 ;
        RECT 0.37 0.402 0.398 0.43 ;
        RECT 0.462 0.466 0.49 0.494 ;
        RECT 0.626 0.402 0.654 0.43 ;
        RECT 0.762 0.402 0.79 0.43 ;
        RECT 0.946 0.402 0.974 0.43 ;
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.238 0.13 ;
        RECT 0.242 0.264 0.27 0.541 ;
        RECT 0.37 0.242 0.398 0.502 ;
        RECT 0.462 0.372 0.494 0.51 ;
        RECT 0.626 0.166 0.654 0.194 ;
        RECT 0.626 0.194 0.654 0.556 ;
        RECT 0.626 0.556 0.654 0.592 ;
        RECT 0.654 0.166 0.75 0.194 ;
        RECT 0.654 0.556 0.75 0.592 ;
        RECT 0.75 0.166 0.755 0.194 ;
        RECT 0.754 0.248 0.79 0.463 ;
        RECT 0.754 0.463 0.79 0.502 ;
        RECT 0.79 0.463 0.8179 0.502 ;
        RECT 0.8179 0.463 0.846 0.502 ;
        RECT 0.8179 0.502 0.846 0.584 ;
        RECT 0.946 0.226 0.974 0.574 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.628 ;
        RECT 0.178 0.628 0.206 0.676 ;
        RECT 0.206 0.166 0.302 0.194 ;
        RECT 0.206 0.628 0.302 0.676 ;
        RECT 0.302 0.628 0.366 0.676 ;
        RECT 0.306 0.307 0.334 0.546 ;
        RECT 0.306 0.546 0.334 0.574 ;
        RECT 0.334 0.546 0.558 0.574 ;
        RECT 0.558 0.184 0.59 0.307 ;
        RECT 0.558 0.307 0.59 0.546 ;
        RECT 0.558 0.546 0.59 0.574 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.334 ;
        RECT 0.462 0.1019 0.466 0.13 ;
        RECT 0.466 0.1019 0.882 0.13 ;
        RECT 0.466 0.628 0.882 0.676 ;
        RECT 0.882 0.1019 0.91 0.13 ;
        RECT 0.882 0.13 0.91 0.334 ;
        RECT 0.882 0.334 0.91 0.628 ;
        RECT 0.882 0.628 0.91 0.676 ;
  END
END CLKGATETST_X1_12T

MACRO DFFRNQ_X1_12T
  CLASS core ;
  FOREIGN DFFRNQ_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.496 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.704 0.274 1.1339 0.302 ;
        RECT 1.1339 0.274 1.326 0.302 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.064 1.616 0.704 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.8139 0.796 ;
        RECT 0.8139 0.74 0.91 0.796 ;
        RECT 0.91 0.74 0.974 0.796 ;
        RECT 0.974 0.74 1.102 0.796 ;
        RECT 1.102 0.74 1.188 0.796 ;
        RECT 1.188 0.74 1.488 0.796 ;
        RECT 1.488 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.21 1.1339 0.238 ;
        RECT 0.082 0.53 1.1339 0.558 ;
      LAYER MINT1 ;
        RECT 0.146 0.21 1.1339 0.238 ;
        RECT 0.082 0.53 1.1339 0.558 ;
      LAYER M1 ;
        RECT 0.178 0.072 0.206 0.6959 ;
        RECT 0.306 0.072 0.334 0.6959 ;
        RECT 0.53 0.623 0.8139 0.681 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.438 ;
        RECT 0.434 0.438 0.462 0.67 ;
        RECT 0.462 0.1019 0.8 0.13 ;
        RECT 0.8 0.1019 0.828 0.13 ;
        RECT 0.8 0.13 0.828 0.438 ;
        RECT 0.576 0.33 0.604 0.506 ;
        RECT 0.576 0.506 0.604 0.534 ;
        RECT 0.604 0.506 0.882 0.534 ;
        RECT 0.882 0.072 0.91 0.33 ;
        RECT 0.882 0.33 0.91 0.506 ;
        RECT 0.882 0.506 0.91 0.534 ;
        RECT 0.882 0.534 0.91 0.672 ;
        RECT 1.01 0.1019 1.038 0.13 ;
        RECT 1.01 0.13 1.038 0.366 ;
        RECT 1.01 0.366 1.038 0.67 ;
        RECT 1.038 0.1019 1.335 0.13 ;
        RECT 1.335 0.1019 1.363 0.13 ;
        RECT 1.335 0.13 1.363 0.366 ;
        RECT 1.224 0.394 1.252 0.638 ;
        RECT 1.224 0.638 1.252 0.666 ;
        RECT 1.252 0.638 1.458 0.666 ;
        RECT 1.458 0.072 1.486 0.132 ;
        RECT 1.458 0.132 1.486 0.394 ;
        RECT 1.458 0.394 1.486 0.638 ;
        RECT 1.458 0.638 1.486 0.666 ;
        RECT 1.486 0.132 1.488 0.394 ;
        RECT 1.486 0.394 1.488 0.638 ;
        RECT 1.486 0.638 1.488 0.666 ;
        RECT 0.048 0.085 0.08 0.1409 ;
        RECT 0.048 0.1409 0.08 0.169 ;
        RECT 0.048 0.5669 0.08 0.606 ;
        RECT 0.048 0.606 0.08 0.686 ;
        RECT 0.08 0.1409 0.114 0.169 ;
        RECT 0.08 0.5669 0.114 0.606 ;
        RECT 0.114 0.1409 0.1419 0.169 ;
        RECT 0.114 0.169 0.1419 0.5669 ;
        RECT 0.114 0.5669 0.1419 0.606 ;
        RECT 0.37 0.194 0.398 0.494 ;
        RECT 0.498 0.402 0.526 0.574 ;
        RECT 0.526 0.194 0.558 0.294 ;
        RECT 0.736 0.258 0.764 0.438 ;
        RECT 0.946 0.274 0.974 0.578 ;
        RECT 1.074 0.1739 1.102 0.317 ;
        RECT 1.074 0.46 1.102 0.622 ;
        RECT 1.156 0.166 1.188 0.686 ;
        RECT 1.266 0.1739 1.294 0.318 ;
      LAYER V1 ;
        RECT 0.114 0.53 0.1419 0.558 ;
        RECT 0.178 0.21 0.206 0.238 ;
        RECT 0.37 0.21 0.398 0.238 ;
        RECT 0.498 0.53 0.526 0.558 ;
        RECT 0.53 0.21 0.558 0.238 ;
        RECT 0.736 0.274 0.764 0.302 ;
        RECT 0.946 0.53 0.974 0.558 ;
        RECT 1.074 0.21 1.102 0.238 ;
        RECT 1.074 0.53 1.102 0.558 ;
        RECT 1.266 0.274 1.294 0.302 ;
      LAYER M1 ;
        RECT 0.178 0.072 0.206 0.6959 ;
        RECT 0.306 0.072 0.334 0.6959 ;
        RECT 0.53 0.623 0.8139 0.681 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.438 ;
        RECT 0.434 0.438 0.462 0.67 ;
        RECT 0.462 0.1019 0.8 0.13 ;
        RECT 0.8 0.1019 0.828 0.13 ;
        RECT 0.8 0.13 0.828 0.438 ;
        RECT 0.576 0.33 0.604 0.506 ;
        RECT 0.576 0.506 0.604 0.534 ;
        RECT 0.604 0.506 0.882 0.534 ;
        RECT 0.882 0.072 0.91 0.33 ;
        RECT 0.882 0.33 0.91 0.506 ;
        RECT 0.882 0.506 0.91 0.534 ;
        RECT 0.882 0.534 0.91 0.672 ;
        RECT 1.01 0.1019 1.038 0.13 ;
        RECT 1.01 0.13 1.038 0.366 ;
        RECT 1.01 0.366 1.038 0.67 ;
        RECT 1.038 0.1019 1.335 0.13 ;
        RECT 1.335 0.1019 1.363 0.13 ;
        RECT 1.335 0.13 1.363 0.366 ;
        RECT 1.224 0.394 1.252 0.638 ;
        RECT 1.224 0.638 1.252 0.666 ;
        RECT 1.252 0.638 1.458 0.666 ;
        RECT 1.458 0.072 1.486 0.132 ;
        RECT 1.458 0.132 1.486 0.394 ;
        RECT 1.458 0.394 1.486 0.638 ;
        RECT 1.458 0.638 1.486 0.666 ;
        RECT 1.486 0.132 1.488 0.394 ;
        RECT 1.486 0.394 1.488 0.638 ;
        RECT 1.486 0.638 1.488 0.666 ;
        RECT 0.048 0.085 0.08 0.1409 ;
        RECT 0.048 0.1409 0.08 0.169 ;
        RECT 0.048 0.5669 0.08 0.606 ;
        RECT 0.048 0.606 0.08 0.686 ;
        RECT 0.08 0.1409 0.114 0.169 ;
        RECT 0.08 0.5669 0.114 0.606 ;
        RECT 0.114 0.1409 0.1419 0.169 ;
        RECT 0.114 0.169 0.1419 0.5669 ;
        RECT 0.114 0.5669 0.1419 0.606 ;
        RECT 0.37 0.194 0.398 0.494 ;
        RECT 0.498 0.402 0.526 0.574 ;
        RECT 0.526 0.194 0.558 0.294 ;
        RECT 0.736 0.258 0.764 0.438 ;
        RECT 0.946 0.274 0.974 0.578 ;
        RECT 1.074 0.1739 1.102 0.317 ;
        RECT 1.074 0.46 1.102 0.622 ;
        RECT 1.156 0.166 1.188 0.686 ;
        RECT 1.266 0.1739 1.294 0.318 ;
  END
END DFFRNQ_X1_12T

MACRO DFFSNQ_X1_12T
  CLASS core ;
  FOREIGN DFFSNQ_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.496 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.722 0.274 1.1339 0.302 ;
        RECT 1.1339 0.274 1.326 0.302 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.064 1.616 0.704 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.554 0.796 ;
        RECT 0.554 0.74 0.91 0.796 ;
        RECT 0.91 0.74 0.974 0.796 ;
        RECT 0.974 0.74 1.106 0.796 ;
        RECT 1.106 0.74 1.3899 0.796 ;
        RECT 1.3899 0.74 1.488 0.796 ;
        RECT 1.488 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.21 1.1339 0.238 ;
        RECT 0.082 0.53 1.1339 0.558 ;
      LAYER MINT1 ;
        RECT 0.146 0.21 1.1339 0.238 ;
        RECT 0.082 0.53 1.1339 0.558 ;
      LAYER M1 ;
        RECT 0.178 0.072 0.206 0.6959 ;
        RECT 0.306 0.072 0.334 0.6959 ;
        RECT 0.434 0.122 0.462 0.15 ;
        RECT 0.434 0.15 0.462 0.366 ;
        RECT 0.434 0.366 0.462 0.67 ;
        RECT 0.462 0.122 0.8179 0.15 ;
        RECT 0.8179 0.122 0.846 0.15 ;
        RECT 0.8179 0.15 0.846 0.366 ;
        RECT 0.946 0.274 0.974 0.574 ;
        RECT 1.074 0.194 1.106 0.325 ;
        RECT 1.074 0.393 1.106 0.594 ;
        RECT 1.266 0.186 1.294 0.318 ;
        RECT 1.202 0.394 1.23 0.574 ;
        RECT 1.202 0.574 1.23 0.602 ;
        RECT 1.23 0.574 1.458 0.602 ;
        RECT 1.458 0.072 1.486 0.132 ;
        RECT 1.458 0.132 1.486 0.394 ;
        RECT 1.458 0.394 1.486 0.574 ;
        RECT 1.458 0.574 1.486 0.602 ;
        RECT 1.486 0.132 1.488 0.394 ;
        RECT 1.486 0.394 1.488 0.574 ;
        RECT 1.486 0.574 1.488 0.602 ;
        RECT 0.045 0.082 0.048 0.138 ;
        RECT 0.045 0.138 0.048 0.177 ;
        RECT 0.048 0.082 0.08 0.138 ;
        RECT 0.048 0.138 0.08 0.177 ;
        RECT 0.048 0.5669 0.08 0.606 ;
        RECT 0.048 0.606 0.08 0.686 ;
        RECT 0.08 0.082 0.083 0.138 ;
        RECT 0.08 0.138 0.083 0.177 ;
        RECT 0.08 0.5669 0.083 0.606 ;
        RECT 0.083 0.138 0.114 0.177 ;
        RECT 0.083 0.5669 0.114 0.606 ;
        RECT 0.114 0.138 0.1419 0.177 ;
        RECT 0.114 0.177 0.1419 0.5669 ;
        RECT 0.114 0.5669 0.1419 0.606 ;
        RECT 0.37 0.194 0.398 0.494 ;
        RECT 0.498 0.402 0.526 0.59 ;
        RECT 0.526 0.194 0.554 0.305 ;
        RECT 0.754 0.258 0.782 0.366 ;
        RECT 0.608 0.274 0.636 0.574 ;
        RECT 0.608 0.574 0.636 0.602 ;
        RECT 0.636 0.574 0.878 0.602 ;
        RECT 0.878 0.574 0.882 0.602 ;
        RECT 0.878 0.602 0.882 0.686 ;
        RECT 0.882 0.096 0.91 0.274 ;
        RECT 0.882 0.274 0.91 0.574 ;
        RECT 0.882 0.574 0.91 0.602 ;
        RECT 0.882 0.602 0.91 0.686 ;
        RECT 1.01 0.114 1.038 0.1419 ;
        RECT 1.01 0.1419 1.038 0.366 ;
        RECT 1.01 0.366 1.038 0.672 ;
        RECT 1.038 0.114 1.352 0.1419 ;
        RECT 1.352 0.114 1.3799 0.1419 ;
        RECT 1.352 0.1419 1.3799 0.366 ;
        RECT 1.106 0.638 1.3899 0.666 ;
      LAYER V1 ;
        RECT 0.114 0.53 0.1419 0.558 ;
        RECT 0.178 0.21 0.206 0.238 ;
        RECT 0.37 0.21 0.398 0.238 ;
        RECT 0.498 0.53 0.526 0.558 ;
        RECT 0.526 0.21 0.554 0.238 ;
        RECT 0.754 0.274 0.782 0.302 ;
        RECT 0.946 0.53 0.974 0.558 ;
        RECT 1.074 0.21 1.102 0.238 ;
        RECT 1.074 0.53 1.102 0.558 ;
        RECT 1.266 0.274 1.294 0.302 ;
      LAYER M1 ;
        RECT 0.178 0.072 0.206 0.6959 ;
        RECT 0.306 0.072 0.334 0.6959 ;
        RECT 0.434 0.122 0.462 0.15 ;
        RECT 0.434 0.15 0.462 0.366 ;
        RECT 0.434 0.366 0.462 0.67 ;
        RECT 0.462 0.122 0.8179 0.15 ;
        RECT 0.8179 0.122 0.846 0.15 ;
        RECT 0.8179 0.15 0.846 0.366 ;
        RECT 0.946 0.274 0.974 0.574 ;
        RECT 1.074 0.194 1.106 0.325 ;
        RECT 1.074 0.393 1.106 0.594 ;
        RECT 1.266 0.186 1.294 0.318 ;
        RECT 1.202 0.394 1.23 0.574 ;
        RECT 1.202 0.574 1.23 0.602 ;
        RECT 1.23 0.574 1.458 0.602 ;
        RECT 1.458 0.072 1.486 0.132 ;
        RECT 1.458 0.132 1.486 0.394 ;
        RECT 1.458 0.394 1.486 0.574 ;
        RECT 1.458 0.574 1.486 0.602 ;
        RECT 1.486 0.132 1.488 0.394 ;
        RECT 1.486 0.394 1.488 0.574 ;
        RECT 1.486 0.574 1.488 0.602 ;
        RECT 0.045 0.082 0.048 0.138 ;
        RECT 0.045 0.138 0.048 0.177 ;
        RECT 0.048 0.082 0.08 0.138 ;
        RECT 0.048 0.138 0.08 0.177 ;
        RECT 0.048 0.5669 0.08 0.606 ;
        RECT 0.048 0.606 0.08 0.686 ;
        RECT 0.08 0.082 0.083 0.138 ;
        RECT 0.08 0.138 0.083 0.177 ;
        RECT 0.08 0.5669 0.083 0.606 ;
        RECT 0.083 0.138 0.114 0.177 ;
        RECT 0.083 0.5669 0.114 0.606 ;
        RECT 0.114 0.138 0.1419 0.177 ;
        RECT 0.114 0.177 0.1419 0.5669 ;
        RECT 0.114 0.5669 0.1419 0.606 ;
        RECT 0.37 0.194 0.398 0.494 ;
        RECT 0.498 0.402 0.526 0.59 ;
        RECT 0.526 0.194 0.554 0.305 ;
        RECT 0.754 0.258 0.782 0.366 ;
        RECT 0.608 0.274 0.636 0.574 ;
        RECT 0.608 0.574 0.636 0.602 ;
        RECT 0.636 0.574 0.878 0.602 ;
        RECT 0.878 0.574 0.882 0.602 ;
        RECT 0.878 0.602 0.882 0.686 ;
        RECT 0.882 0.096 0.91 0.274 ;
        RECT 0.882 0.274 0.91 0.574 ;
        RECT 0.882 0.574 0.91 0.602 ;
        RECT 0.882 0.602 0.91 0.686 ;
        RECT 1.01 0.114 1.038 0.1419 ;
        RECT 1.01 0.1419 1.038 0.366 ;
        RECT 1.01 0.366 1.038 0.672 ;
        RECT 1.038 0.114 1.352 0.1419 ;
        RECT 1.352 0.114 1.3799 0.1419 ;
        RECT 1.352 0.1419 1.3799 0.366 ;
        RECT 1.106 0.638 1.3899 0.666 ;
  END
END DFFSNQ_X1_12T

MACRO FA_X1_12T
  CLASS core ;
  FOREIGN FA_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.304 BY 0.512 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.21 0.466 1.098 0.494 ;
      LAYER V1 ;
        RECT 0.656 0.466 0.684 0.494 ;
        RECT 1.038 0.466 1.066 0.494 ;
      LAYER M1 ;
        RECT 0.656 0.402 0.684 0.526 ;
        RECT 1.038 0.274 1.074 0.526 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.274 0.274 0.789 0.302 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.146 0.21 1.262 0.238 ;
      LAYER V1 ;
        RECT 0.178 0.21 0.206 0.238 ;
        RECT 0.58 0.21 0.608 0.238 ;
        RECT 1.202 0.21 1.23 0.238 ;
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.59 ;
        RECT 0.58 0.194 0.608 0.366 ;
        RECT 1.202 0.178 1.23 0.366 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.458 0.114 1.486 0.654 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8179 0.207 0.846 0.64 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.656 0.796 ;
        RECT 0.656 0.74 0.767 0.796 ;
        RECT 0.767 0.74 1.038 0.796 ;
        RECT 1.038 0.74 1.084 0.796 ;
        RECT 1.084 0.74 1.166 0.796 ;
        RECT 1.166 0.74 1.289 0.796 ;
        RECT 1.289 0.74 1.358 0.796 ;
        RECT 1.358 0.74 1.546 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.546 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.082 0.402 1.321 0.43 ;
        RECT 0.402 0.338 1.3899 0.366 ;
      LAYER MINT1 ;
        RECT 0.082 0.402 1.321 0.43 ;
        RECT 0.402 0.338 1.3899 0.366 ;
      LAYER M1 ;
        RECT 0.027 0.178 0.065 0.338 ;
        RECT 0.027 0.338 0.065 0.366 ;
        RECT 0.065 0.338 0.103 0.366 ;
        RECT 0.103 0.338 0.1419 0.366 ;
        RECT 0.103 0.366 0.1419 0.462 ;
        RECT 0.242 0.274 0.27 0.59 ;
        RECT 0.424 0.274 0.462 0.507 ;
        RECT 0.37 0.097 0.618 0.135 ;
        RECT 0.37 0.575 0.402 0.603 ;
        RECT 0.37 0.603 0.402 0.6979 ;
        RECT 0.402 0.575 0.624 0.603 ;
        RECT 0.624 0.575 0.656 0.603 ;
        RECT 0.624 0.603 0.656 0.6979 ;
        RECT 0.624 0.6979 0.656 0.704 ;
        RECT 0.729 0.244 0.767 0.464 ;
        RECT 0.882 0.194 0.91 0.366 ;
        RECT 0.882 0.562 0.91 0.59 ;
        RECT 0.882 0.59 0.91 0.6959 ;
        RECT 0.91 0.562 1.01 0.59 ;
        RECT 1.01 0.562 1.038 0.59 ;
        RECT 1.01 0.59 1.038 0.6959 ;
        RECT 1.1379 0.072 1.166 0.6959 ;
        RECT 1.2609 0.386 1.289 0.59 ;
        RECT 0.306 0.096 0.334 0.672 ;
        RECT 0.498 0.274 0.526 0.507 ;
        RECT 0.946 0.274 0.984 0.494 ;
        RECT 0.846 0.1 1.084 0.132 ;
        RECT 1.33 0.274 1.358 0.526 ;
      LAYER V1 ;
        RECT 0.114 0.402 0.1419 0.43 ;
        RECT 0.242 0.466 0.27 0.494 ;
        RECT 0.306 0.274 0.334 0.302 ;
        RECT 0.434 0.338 0.462 0.366 ;
        RECT 0.498 0.402 0.526 0.43 ;
        RECT 0.729 0.274 0.757 0.302 ;
        RECT 0.882 0.21 0.91 0.238 ;
        RECT 0.956 0.402 0.984 0.43 ;
        RECT 1.1379 0.338 1.166 0.366 ;
        RECT 1.2609 0.402 1.289 0.43 ;
        RECT 1.33 0.338 1.358 0.366 ;
      LAYER M1 ;
        RECT 0.027 0.178 0.065 0.338 ;
        RECT 0.027 0.338 0.065 0.366 ;
        RECT 0.065 0.338 0.103 0.366 ;
        RECT 0.103 0.338 0.1419 0.366 ;
        RECT 0.103 0.366 0.1419 0.462 ;
        RECT 0.242 0.274 0.27 0.59 ;
        RECT 0.424 0.274 0.462 0.507 ;
        RECT 0.37 0.097 0.618 0.135 ;
        RECT 0.37 0.575 0.402 0.603 ;
        RECT 0.37 0.603 0.402 0.6979 ;
        RECT 0.402 0.575 0.624 0.603 ;
        RECT 0.624 0.575 0.656 0.603 ;
        RECT 0.624 0.603 0.656 0.6979 ;
        RECT 0.624 0.6979 0.656 0.704 ;
        RECT 0.729 0.244 0.767 0.464 ;
        RECT 0.882 0.194 0.91 0.366 ;
        RECT 0.882 0.562 0.91 0.59 ;
        RECT 0.882 0.59 0.91 0.6959 ;
        RECT 0.91 0.562 1.01 0.59 ;
        RECT 1.01 0.562 1.038 0.59 ;
        RECT 1.01 0.59 1.038 0.6959 ;
        RECT 1.1379 0.072 1.166 0.6959 ;
        RECT 1.2609 0.386 1.289 0.59 ;
        RECT 0.306 0.096 0.334 0.672 ;
        RECT 0.498 0.274 0.526 0.507 ;
        RECT 0.946 0.274 0.984 0.494 ;
        RECT 0.846 0.1 1.084 0.132 ;
        RECT 1.33 0.274 1.358 0.526 ;
  END
END FA_X1_12T

MACRO FILLTIE_12T
  CLASS core ;
  FOREIGN FILLTIE_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.867 BY 0.512 ;
  OBS
      LAYER M1 ;
        RECT -0.01 -0.028 0.588 0.028 ;
        RECT -0.01 0.74 0.588 0.796 ;
      LAYER M1 ;
        RECT -0.01 -0.028 0.588 0.028 ;
        RECT -0.01 0.74 0.588 0.796 ;
  END
END FILLTIE_12T

MACRO FILL_X1_12T
  CLASS core ;
  FOREIGN FILL_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.138 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.138 0.028 ;
    END
  END VSS
END FILL_X1_12T

MACRO FILL_X2_12T
  CLASS core ;
  FOREIGN FILL_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.288 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
END FILL_X2_12T

MACRO FILL_X4_12T
  CLASS core ;
  FOREIGN FILL_X4_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.48 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
END FILL_X4_12T

MACRO FILL_X8_12T
  CLASS core ;
  FOREIGN FILL_X8_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
END FILL_X8_12T

MACRO FILL_X16_12T
  CLASS core ;
  FOREIGN FILL_X16_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.632 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.098 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.098 0.028 ;
    END
  END VSS
END FILL_X16_12T

MACRO HA_X1_12T
  CLASS core ;
  FOREIGN HA_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.248 BY 0.512 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.274 0.27 0.556 ;
        RECT 0.242 0.556 0.27 0.584 ;
        RECT 0.27 0.556 0.434 0.584 ;
        RECT 0.434 0.274 0.462 0.556 ;
        RECT 0.434 0.556 0.462 0.584 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.512 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.082 0.078 0.638 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.754 0.18 0.782 0.638 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.596 0.796 ;
        RECT 0.596 0.74 0.66 0.796 ;
        RECT 0.66 0.74 0.842 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.842 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.338 0.1019 0.622 0.13 ;
        RECT 0.406 0.184 0.498 0.216 ;
        RECT 0.498 0.184 0.53 0.216 ;
        RECT 0.498 0.216 0.53 0.462 ;
        RECT 0.498 0.462 0.53 0.602 ;
        RECT 0.53 0.184 0.632 0.216 ;
        RECT 0.632 0.184 0.66 0.216 ;
        RECT 0.632 0.216 0.66 0.462 ;
        RECT 0.114 0.166 0.1419 0.198 ;
        RECT 0.114 0.198 0.1419 0.274 ;
        RECT 0.114 0.274 0.1419 0.638 ;
        RECT 0.114 0.638 0.1419 0.666 ;
        RECT 0.1419 0.166 0.37 0.198 ;
        RECT 0.1419 0.638 0.37 0.666 ;
        RECT 0.37 0.638 0.5659 0.666 ;
        RECT 0.5659 0.274 0.596 0.638 ;
        RECT 0.5659 0.638 0.596 0.666 ;
      LAYER M1 ;
        RECT 0.338 0.1019 0.622 0.13 ;
        RECT 0.406 0.184 0.498 0.216 ;
        RECT 0.498 0.184 0.53 0.216 ;
        RECT 0.498 0.216 0.53 0.462 ;
        RECT 0.498 0.462 0.53 0.602 ;
        RECT 0.53 0.184 0.632 0.216 ;
        RECT 0.632 0.184 0.66 0.216 ;
        RECT 0.632 0.216 0.66 0.462 ;
        RECT 0.114 0.166 0.1419 0.198 ;
        RECT 0.114 0.198 0.1419 0.274 ;
        RECT 0.114 0.274 0.1419 0.638 ;
        RECT 0.114 0.638 0.1419 0.666 ;
        RECT 0.1419 0.166 0.37 0.198 ;
        RECT 0.1419 0.638 0.37 0.666 ;
        RECT 0.37 0.638 0.5659 0.666 ;
        RECT 0.5659 0.274 0.596 0.638 ;
        RECT 0.5659 0.638 0.596 0.666 ;
  END
END HA_X1_12T

MACRO INV_X1_12T
  CLASS core ;
  FOREIGN INV_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.288 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.114 0.1419 0.64 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
END INV_X1_12T

MACRO INV_X2_12T
  CLASS core ;
  FOREIGN INV_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.13 0.1419 0.576 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
END INV_X2_12T

MACRO INV_X4_12T
  CLASS core ;
  FOREIGN INV_X4_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.256 0.08 0.368 ;
        RECT 0.048 0.368 0.08 0.396 ;
        RECT 0.048 0.396 0.08 0.512 ;
        RECT 0.08 0.368 0.238 0.396 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.1419 0.059 0.2 ;
        RECT 0.059 0.1419 0.306 0.2 ;
        RECT 0.059 0.5679 0.306 0.626 ;
        RECT 0.306 0.1419 0.334 0.2 ;
        RECT 0.306 0.2 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.626 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END INV_X4_12T

MACRO INV_X8_12T
  CLASS core ;
  FOREIGN INV_X8_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.96 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.194 0.1419 0.396 ;
        RECT 0.114 0.396 0.1419 0.455 ;
        RECT 0.114 0.455 0.1419 0.576 ;
        RECT 0.1419 0.396 0.462 0.455 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.631 0.054 0.659 ;
        RECT 0.054 0.11 0.557 0.138 ;
        RECT 0.054 0.631 0.557 0.659 ;
        RECT 0.557 0.11 0.595 0.138 ;
        RECT 0.557 0.138 0.595 0.631 ;
        RECT 0.557 0.631 0.595 0.659 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
END INV_X8_12T

MACRO INV_X12_12T
  CLASS core ;
  FOREIGN INV_X12_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.344 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.1419 0.368 ;
        RECT 0.114 0.368 0.1419 0.396 ;
        RECT 0.114 0.396 0.1419 0.576 ;
        RECT 0.1419 0.368 0.686 0.396 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.1019 0.8129 0.13 ;
        RECT 0.054 0.636 0.8129 0.668 ;
        RECT 0.8129 0.1019 0.851 0.13 ;
        RECT 0.8129 0.13 0.851 0.636 ;
        RECT 0.8129 0.636 0.851 0.668 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
END INV_X12_12T

MACRO LHQ_X1_12T
  CLASS core ;
  FOREIGN LHQ_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.344 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.16 0.27 0.512 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8179 0.13 0.846 0.638 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.782 0.796 ;
        RECT 0.782 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.556 0.05 0.584 ;
        RECT 0.048 0.584 0.05 0.704 ;
        RECT 0.05 0.064 0.078 0.092 ;
        RECT 0.05 0.092 0.078 0.184 ;
        RECT 0.05 0.184 0.078 0.212 ;
        RECT 0.05 0.556 0.078 0.584 ;
        RECT 0.05 0.584 0.078 0.704 ;
        RECT 0.078 0.064 0.08 0.092 ;
        RECT 0.078 0.184 0.08 0.212 ;
        RECT 0.078 0.556 0.08 0.584 ;
        RECT 0.078 0.584 0.08 0.704 ;
        RECT 0.08 0.064 0.114 0.092 ;
        RECT 0.08 0.184 0.114 0.212 ;
        RECT 0.08 0.556 0.114 0.584 ;
        RECT 0.114 0.064 0.1419 0.092 ;
        RECT 0.114 0.184 0.1419 0.212 ;
        RECT 0.114 0.212 0.1419 0.322 ;
        RECT 0.114 0.322 0.1419 0.35 ;
        RECT 0.114 0.35 0.1419 0.414 ;
        RECT 0.114 0.414 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.064 0.324 0.092 ;
        RECT 0.324 0.064 0.352 0.092 ;
        RECT 0.324 0.092 0.352 0.184 ;
        RECT 0.324 0.184 0.352 0.212 ;
        RECT 0.324 0.212 0.352 0.322 ;
        RECT 0.324 0.322 0.352 0.35 ;
        RECT 0.352 0.322 0.37 0.35 ;
        RECT 0.37 0.322 0.398 0.35 ;
        RECT 0.37 0.35 0.398 0.414 ;
        RECT 0.53 0.114 0.558 0.1419 ;
        RECT 0.53 0.1419 0.558 0.494 ;
        RECT 0.558 0.114 0.6899 0.1419 ;
        RECT 0.6899 0.114 0.718 0.1419 ;
        RECT 0.6899 0.1419 0.718 0.494 ;
        RECT 0.6899 0.494 0.718 0.593 ;
        RECT 0.178 0.136 0.206 0.46 ;
        RECT 0.178 0.46 0.206 0.556 ;
        RECT 0.178 0.556 0.206 0.584 ;
        RECT 0.206 0.556 0.306 0.584 ;
        RECT 0.306 0.46 0.34 0.556 ;
        RECT 0.306 0.556 0.34 0.584 ;
        RECT 0.274 0.638 0.388 0.666 ;
        RECT 0.388 0.114 0.466 0.1729 ;
        RECT 0.388 0.638 0.466 0.666 ;
        RECT 0.466 0.114 0.494 0.1729 ;
        RECT 0.466 0.1729 0.494 0.306 ;
        RECT 0.466 0.306 0.494 0.637 ;
        RECT 0.466 0.637 0.494 0.638 ;
        RECT 0.466 0.638 0.494 0.666 ;
        RECT 0.494 0.637 0.754 0.638 ;
        RECT 0.494 0.638 0.754 0.666 ;
        RECT 0.754 0.306 0.782 0.637 ;
        RECT 0.754 0.637 0.782 0.638 ;
        RECT 0.754 0.638 0.782 0.666 ;
      LAYER M1 ;
        RECT 0.048 0.556 0.05 0.584 ;
        RECT 0.048 0.584 0.05 0.704 ;
        RECT 0.05 0.064 0.078 0.092 ;
        RECT 0.05 0.092 0.078 0.184 ;
        RECT 0.05 0.184 0.078 0.212 ;
        RECT 0.05 0.556 0.078 0.584 ;
        RECT 0.05 0.584 0.078 0.704 ;
        RECT 0.078 0.064 0.08 0.092 ;
        RECT 0.078 0.184 0.08 0.212 ;
        RECT 0.078 0.556 0.08 0.584 ;
        RECT 0.078 0.584 0.08 0.704 ;
        RECT 0.08 0.064 0.114 0.092 ;
        RECT 0.08 0.184 0.114 0.212 ;
        RECT 0.08 0.556 0.114 0.584 ;
        RECT 0.114 0.064 0.1419 0.092 ;
        RECT 0.114 0.184 0.1419 0.212 ;
        RECT 0.114 0.212 0.1419 0.322 ;
        RECT 0.114 0.322 0.1419 0.35 ;
        RECT 0.114 0.35 0.1419 0.414 ;
        RECT 0.114 0.414 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.064 0.324 0.092 ;
        RECT 0.324 0.064 0.352 0.092 ;
        RECT 0.324 0.092 0.352 0.184 ;
        RECT 0.324 0.184 0.352 0.212 ;
        RECT 0.324 0.212 0.352 0.322 ;
        RECT 0.324 0.322 0.352 0.35 ;
        RECT 0.352 0.322 0.37 0.35 ;
        RECT 0.37 0.322 0.398 0.35 ;
        RECT 0.37 0.35 0.398 0.414 ;
        RECT 0.53 0.114 0.558 0.1419 ;
        RECT 0.53 0.1419 0.558 0.494 ;
        RECT 0.558 0.114 0.6899 0.1419 ;
        RECT 0.6899 0.114 0.718 0.1419 ;
        RECT 0.6899 0.1419 0.718 0.494 ;
        RECT 0.6899 0.494 0.718 0.593 ;
        RECT 0.178 0.136 0.206 0.46 ;
        RECT 0.178 0.46 0.206 0.556 ;
        RECT 0.178 0.556 0.206 0.584 ;
        RECT 0.206 0.556 0.306 0.584 ;
        RECT 0.306 0.46 0.34 0.556 ;
        RECT 0.306 0.556 0.34 0.584 ;
        RECT 0.274 0.638 0.388 0.666 ;
        RECT 0.388 0.114 0.466 0.1729 ;
        RECT 0.388 0.638 0.466 0.666 ;
        RECT 0.466 0.114 0.494 0.1729 ;
        RECT 0.466 0.1729 0.494 0.306 ;
        RECT 0.466 0.306 0.494 0.637 ;
        RECT 0.466 0.637 0.494 0.638 ;
        RECT 0.466 0.638 0.494 0.666 ;
        RECT 0.494 0.637 0.754 0.638 ;
        RECT 0.494 0.638 0.754 0.666 ;
        RECT 0.754 0.306 0.782 0.637 ;
        RECT 0.754 0.637 0.782 0.638 ;
        RECT 0.754 0.638 0.782 0.666 ;
  END
END LHQ_X1_12T

MACRO MUX2_X1_12T
  CLASS core ;
  FOREIGN MUX2_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.248 BY 0.512 ;
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.242 0.59 0.526 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.448 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.118 0.658 0.394 0.686 ;
      LAYER V1 ;
        RECT 0.15 0.658 0.206 0.686 ;
      LAYER M1 ;
        RECT 0.027 0.242 0.055 0.658 ;
        RECT 0.027 0.658 0.055 0.686 ;
        RECT 0.055 0.658 0.222 0.686 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.6899 0.192 0.718 0.638 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.462 0.796 ;
        RECT 0.462 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.782 0.796 ;
        RECT 0.782 0.74 0.842 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.842 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.274 0.338 0.558 0.366 ;
      LAYER MINT1 ;
        RECT 0.274 0.338 0.558 0.366 ;
      LAYER M1 ;
        RECT 0.08 0.162 0.099 0.19 ;
        RECT 0.099 0.162 0.157 0.19 ;
        RECT 0.099 0.492 0.157 0.52 ;
        RECT 0.099 0.52 0.157 0.576 ;
        RECT 0.157 0.162 0.306 0.19 ;
        RECT 0.157 0.492 0.306 0.52 ;
        RECT 0.306 0.162 0.334 0.19 ;
        RECT 0.306 0.19 0.334 0.492 ;
        RECT 0.306 0.492 0.334 0.52 ;
        RECT 0.29 0.658 0.434 0.704 ;
        RECT 0.434 0.306 0.462 0.658 ;
        RECT 0.434 0.658 0.462 0.704 ;
        RECT 0.498 0.274 0.526 0.428 ;
        RECT 0.37 0.0869 0.398 0.146 ;
        RECT 0.37 0.146 0.398 0.494 ;
        RECT 0.37 0.494 0.398 0.614 ;
        RECT 0.398 0.0869 0.754 0.146 ;
        RECT 0.754 0.0869 0.782 0.146 ;
        RECT 0.754 0.146 0.782 0.494 ;
      LAYER V1 ;
        RECT 0.306 0.338 0.334 0.366 ;
        RECT 0.306 0.658 0.362 0.686 ;
        RECT 0.498 0.338 0.526 0.366 ;
      LAYER M1 ;
        RECT 0.08 0.162 0.099 0.19 ;
        RECT 0.099 0.162 0.157 0.19 ;
        RECT 0.099 0.492 0.157 0.52 ;
        RECT 0.099 0.52 0.157 0.576 ;
        RECT 0.157 0.162 0.306 0.19 ;
        RECT 0.157 0.492 0.306 0.52 ;
        RECT 0.306 0.162 0.334 0.19 ;
        RECT 0.306 0.19 0.334 0.492 ;
        RECT 0.306 0.492 0.334 0.52 ;
        RECT 0.29 0.658 0.434 0.704 ;
        RECT 0.434 0.306 0.462 0.658 ;
        RECT 0.434 0.658 0.462 0.704 ;
        RECT 0.498 0.274 0.526 0.428 ;
        RECT 0.37 0.0869 0.398 0.146 ;
        RECT 0.37 0.146 0.398 0.494 ;
        RECT 0.37 0.494 0.398 0.614 ;
        RECT 0.398 0.0869 0.754 0.146 ;
        RECT 0.754 0.0869 0.782 0.146 ;
        RECT 0.754 0.146 0.782 0.494 ;
  END
END MUX2_X1_12T

MACRO NAND2_X1_12T
  CLASS core ;
  FOREIGN NAND2_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.574 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.574 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.133 0.1419 0.192 ;
        RECT 0.114 0.192 0.1419 0.638 ;
        RECT 0.1419 0.133 0.176 0.192 ;
        RECT 0.176 0.064 0.208 0.133 ;
        RECT 0.176 0.133 0.208 0.192 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
END NAND2_X1_12T

MACRO NAND2_X2_12T
  CLASS core ;
  FOREIGN NAND2_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.225 0.206 0.553 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.274 0.078 0.676 ;
        RECT 0.05 0.676 0.078 0.704 ;
        RECT 0.078 0.676 0.306 0.704 ;
        RECT 0.306 0.274 0.334 0.676 ;
        RECT 0.306 0.676 0.334 0.704 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.123 0.1419 0.181 ;
        RECT 0.114 0.181 0.1419 0.424 ;
        RECT 0.114 0.424 0.1419 0.597 ;
        RECT 0.114 0.597 0.1419 0.64 ;
        RECT 0.1419 0.123 0.242 0.181 ;
        RECT 0.1419 0.597 0.242 0.64 ;
        RECT 0.242 0.123 0.27 0.181 ;
        RECT 0.242 0.424 0.27 0.597 ;
        RECT 0.242 0.597 0.27 0.64 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END NAND2_X2_12T

MACRO NAND3_X1_12T
  CLASS core ;
  FOREIGN NAND3_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.32 0.27 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.255 0.206 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.215 0.078 0.574 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.082 0.1419 0.11 ;
        RECT 0.114 0.11 0.1419 0.256 ;
        RECT 0.114 0.256 0.1419 0.512 ;
        RECT 0.114 0.512 0.1419 0.676 ;
        RECT 0.114 0.676 0.1419 0.704 ;
        RECT 0.1419 0.082 0.242 0.11 ;
        RECT 0.1419 0.676 0.242 0.704 ;
        RECT 0.242 0.064 0.304 0.082 ;
        RECT 0.242 0.082 0.304 0.11 ;
        RECT 0.242 0.676 0.304 0.704 ;
        RECT 0.304 0.064 0.306 0.082 ;
        RECT 0.304 0.082 0.306 0.11 ;
        RECT 0.304 0.11 0.306 0.256 ;
        RECT 0.304 0.676 0.306 0.704 ;
        RECT 0.306 0.064 0.334 0.082 ;
        RECT 0.306 0.082 0.334 0.11 ;
        RECT 0.306 0.11 0.334 0.256 ;
        RECT 0.306 0.512 0.334 0.676 ;
        RECT 0.306 0.676 0.334 0.704 ;
        RECT 0.334 0.064 0.336 0.082 ;
        RECT 0.334 0.082 0.336 0.11 ;
        RECT 0.334 0.11 0.336 0.256 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END NAND3_X1_12T

MACRO NAND3_X2_12T
  CLASS core ;
  FOREIGN NAND3_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.32 0.526 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.301 0.249 0.339 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.512 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.027 0.5679 0.366 0.626 ;
        RECT 0.366 0.5679 0.434 0.626 ;
        RECT 0.434 0.186 0.462 0.5679 ;
        RECT 0.434 0.5679 0.462 0.626 ;
        RECT 0.462 0.5679 0.494 0.626 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.366 0.796 ;
        RECT 0.366 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.111 0.498 0.1409 ;
        RECT 0.498 0.111 0.526 0.1409 ;
        RECT 0.498 0.1409 0.526 0.225 ;
        RECT 0.05 0.177 0.366 0.209 ;
      LAYER M1 ;
        RECT 0.21 0.111 0.498 0.1409 ;
        RECT 0.498 0.111 0.526 0.1409 ;
        RECT 0.498 0.1409 0.526 0.225 ;
        RECT 0.05 0.177 0.366 0.209 ;
  END
END NAND3_X2_12T

MACRO NAND4_X1_12T
  CLASS core ;
  FOREIGN NAND4_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.672 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.256 0.398 0.574 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.448 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.574 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.512 0.1419 0.645 ;
        RECT 0.114 0.645 0.1419 0.704 ;
        RECT 0.1419 0.645 0.306 0.704 ;
        RECT 0.306 0.164 0.334 0.192 ;
        RECT 0.306 0.192 0.334 0.512 ;
        RECT 0.306 0.512 0.334 0.645 ;
        RECT 0.306 0.645 0.334 0.704 ;
        RECT 0.334 0.164 0.365 0.192 ;
        RECT 0.365 0.064 0.403 0.164 ;
        RECT 0.365 0.164 0.403 0.192 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
END NAND4_X1_12T

MACRO NAND4_X2_12T
  CLASS core ;
  FOREIGN NAND4_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.056 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.358 0.594 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.34 0.398 0.526 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.242 0.206 0.512 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.257 0.078 0.512 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.555 0.144 0.576 ;
        RECT 0.112 0.576 0.144 0.638 ;
        RECT 0.112 0.638 0.144 0.666 ;
        RECT 0.144 0.638 0.434 0.666 ;
        RECT 0.434 0.294 0.462 0.322 ;
        RECT 0.434 0.322 0.462 0.548 ;
        RECT 0.434 0.548 0.462 0.555 ;
        RECT 0.434 0.555 0.462 0.576 ;
        RECT 0.434 0.638 0.462 0.666 ;
        RECT 0.462 0.294 0.562 0.322 ;
        RECT 0.462 0.548 0.562 0.555 ;
        RECT 0.462 0.555 0.562 0.576 ;
        RECT 0.462 0.638 0.562 0.666 ;
        RECT 0.562 0.294 0.59 0.322 ;
        RECT 0.562 0.548 0.59 0.555 ;
        RECT 0.562 0.555 0.59 0.576 ;
        RECT 0.562 0.576 0.59 0.638 ;
        RECT 0.562 0.638 0.59 0.666 ;
        RECT 0.59 0.294 0.654 0.322 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.656 0.796 ;
        RECT 0.656 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.43 0.13 ;
        RECT 0.274 0.23 0.624 0.258 ;
        RECT 0.624 0.064 0.656 0.23 ;
        RECT 0.624 0.23 0.656 0.258 ;
        RECT 0.146 0.166 0.494 0.194 ;
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.43 0.13 ;
        RECT 0.274 0.23 0.624 0.258 ;
        RECT 0.624 0.064 0.656 0.23 ;
        RECT 0.624 0.23 0.656 0.258 ;
        RECT 0.146 0.166 0.494 0.194 ;
  END
END NAND4_X2_12T

MACRO NOR2_X1_12T
  CLASS core ;
  FOREIGN NOR2_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.512 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.13 0.1419 0.576 ;
        RECT 0.114 0.576 0.1419 0.635 ;
        RECT 0.1419 0.576 0.176 0.635 ;
        RECT 0.176 0.576 0.208 0.635 ;
        RECT 0.176 0.635 0.208 0.704 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
END NOR2_X1_12T

MACRO NOR2_X2_12T
  CLASS core ;
  FOREIGN NOR2_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.215 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.064 0.078 0.092 ;
        RECT 0.05 0.092 0.078 0.494 ;
        RECT 0.078 0.064 0.306 0.092 ;
        RECT 0.306 0.064 0.334 0.092 ;
        RECT 0.306 0.092 0.334 0.494 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.128 0.1419 0.156 ;
        RECT 0.114 0.156 0.1419 0.3439 ;
        RECT 0.114 0.3439 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.128 0.176 0.156 ;
        RECT 0.1419 0.556 0.176 0.584 ;
        RECT 0.176 0.128 0.208 0.156 ;
        RECT 0.176 0.556 0.208 0.584 ;
        RECT 0.176 0.584 0.208 0.64 ;
        RECT 0.208 0.128 0.242 0.156 ;
        RECT 0.242 0.128 0.27 0.156 ;
        RECT 0.242 0.156 0.27 0.3439 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END NOR2_X2_12T

MACRO NOR3_X1_12T
  CLASS core ;
  FOREIGN NOR3_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.32 0.27 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.553 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.553 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.064 0.1419 0.092 ;
        RECT 0.114 0.092 0.1419 0.256 ;
        RECT 0.114 0.256 0.1419 0.512 ;
        RECT 0.114 0.512 0.1419 0.614 ;
        RECT 0.114 0.614 0.1419 0.642 ;
        RECT 0.1419 0.064 0.303 0.092 ;
        RECT 0.1419 0.614 0.303 0.642 ;
        RECT 0.303 0.064 0.304 0.092 ;
        RECT 0.303 0.092 0.304 0.256 ;
        RECT 0.303 0.614 0.304 0.642 ;
        RECT 0.304 0.064 0.336 0.092 ;
        RECT 0.304 0.092 0.336 0.256 ;
        RECT 0.304 0.512 0.336 0.614 ;
        RECT 0.304 0.614 0.336 0.642 ;
        RECT 0.304 0.642 0.336 0.704 ;
        RECT 0.336 0.064 0.337 0.092 ;
        RECT 0.336 0.092 0.337 0.256 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END NOR3_X1_12T

MACRO NOR3_X2_12T
  CLASS core ;
  FOREIGN NOR3_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.256 0.526 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.513 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.519 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0859 0.154 0.434 0.212 ;
        RECT 0.434 0.154 0.462 0.212 ;
        RECT 0.434 0.212 0.462 0.576 ;
        RECT 0.462 0.154 0.49 0.212 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.627 0.498 0.655 ;
        RECT 0.498 0.516 0.526 0.627 ;
        RECT 0.498 0.627 0.526 0.655 ;
        RECT 0.0859 0.557 0.38 0.591 ;
      LAYER M1 ;
        RECT 0.21 0.627 0.498 0.655 ;
        RECT 0.498 0.516 0.526 0.627 ;
        RECT 0.498 0.627 0.526 0.655 ;
        RECT 0.0859 0.557 0.38 0.591 ;
  END
END NOR3_X2_12T

MACRO NOR4_X1_12T
  CLASS core ;
  FOREIGN NOR4_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.672 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.194 0.398 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.194 0.27 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.574 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.574 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.064 0.1419 0.1019 ;
        RECT 0.114 0.1019 0.1419 0.215 ;
        RECT 0.1419 0.064 0.306 0.1019 ;
        RECT 0.306 0.064 0.334 0.1019 ;
        RECT 0.306 0.1019 0.334 0.215 ;
        RECT 0.306 0.215 0.334 0.576 ;
        RECT 0.306 0.576 0.334 0.604 ;
        RECT 0.334 0.576 0.365 0.604 ;
        RECT 0.365 0.576 0.403 0.604 ;
        RECT 0.365 0.604 0.403 0.704 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
END NOR4_X1_12T

MACRO NOR4_X2_12T
  CLASS core ;
  FOREIGN NOR4_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.056 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.256 0.594 0.406 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.242 0.398 0.438 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.516 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.1019 0.144 0.13 ;
        RECT 0.112 0.13 0.144 0.192 ;
        RECT 0.112 0.192 0.144 0.213 ;
        RECT 0.144 0.1019 0.434 0.13 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.192 0.462 0.213 ;
        RECT 0.434 0.213 0.462 0.22 ;
        RECT 0.434 0.22 0.462 0.442 ;
        RECT 0.434 0.442 0.462 0.47 ;
        RECT 0.462 0.1019 0.562 0.13 ;
        RECT 0.462 0.192 0.562 0.213 ;
        RECT 0.462 0.213 0.562 0.22 ;
        RECT 0.462 0.442 0.562 0.47 ;
        RECT 0.562 0.1019 0.59 0.13 ;
        RECT 0.562 0.13 0.59 0.192 ;
        RECT 0.562 0.192 0.59 0.213 ;
        RECT 0.562 0.213 0.59 0.22 ;
        RECT 0.562 0.442 0.59 0.47 ;
        RECT 0.59 0.442 0.663 0.47 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.43 0.796 ;
        RECT 0.43 0.74 0.494 0.796 ;
        RECT 0.494 0.74 0.656 0.796 ;
        RECT 0.656 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.5699 0.494 0.602 ;
        RECT 0.048 0.555 0.08 0.638 ;
        RECT 0.048 0.638 0.08 0.666 ;
        RECT 0.08 0.638 0.43 0.666 ;
        RECT 0.338 0.506 0.624 0.534 ;
        RECT 0.624 0.506 0.656 0.534 ;
        RECT 0.624 0.534 0.656 0.686 ;
      LAYER M1 ;
        RECT 0.21 0.5699 0.494 0.602 ;
        RECT 0.048 0.555 0.08 0.638 ;
        RECT 0.048 0.638 0.08 0.666 ;
        RECT 0.08 0.638 0.43 0.666 ;
        RECT 0.338 0.506 0.624 0.534 ;
        RECT 0.624 0.506 0.656 0.534 ;
        RECT 0.624 0.534 0.656 0.686 ;
  END
END NOR4_X2_12T

MACRO OAI21_X1_12T
  CLASS core ;
  FOREIGN OAI21_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.634 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.576 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.636 ;
        RECT 0.114 0.636 0.1419 0.668 ;
        RECT 0.1419 0.636 0.298 0.668 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.298 0.796 ;
        RECT 0.298 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.073 0.078 0.155 ;
        RECT 0.05 0.155 0.078 0.187 ;
        RECT 0.078 0.155 0.298 0.187 ;
      LAYER M1 ;
        RECT 0.05 0.073 0.078 0.155 ;
        RECT 0.05 0.155 0.078 0.187 ;
        RECT 0.078 0.155 0.298 0.187 ;
  END
END OAI21_X1_12T

MACRO OAI21_X2_12T
  CLASS core ;
  FOREIGN OAI21_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.365 0.32 0.403 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.2829 ;
        RECT 0.242 0.2829 0.27 0.502 ;
        RECT 0.242 0.502 0.27 0.53 ;
        RECT 0.27 0.502 0.498 0.53 ;
        RECT 0.498 0.2829 0.526 0.502 ;
        RECT 0.498 0.502 0.526 0.53 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.525 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.029 0.5699 0.178 0.602 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.278 ;
        RECT 0.178 0.278 0.206 0.5699 ;
        RECT 0.178 0.5699 0.206 0.602 ;
        RECT 0.206 0.166 0.426 0.194 ;
        RECT 0.206 0.5699 0.426 0.602 ;
        RECT 0.426 0.166 0.434 0.194 ;
        RECT 0.434 0.166 0.462 0.194 ;
        RECT 0.434 0.194 0.462 0.278 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.535 0.796 ;
        RECT 0.535 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.498 0.13 ;
        RECT 0.498 0.1019 0.526 0.13 ;
        RECT 0.498 0.13 0.526 0.213 ;
        RECT 0.498 0.213 0.526 0.215 ;
        RECT 0.146 0.638 0.535 0.666 ;
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.498 0.13 ;
        RECT 0.498 0.1019 0.526 0.13 ;
        RECT 0.498 0.13 0.526 0.213 ;
        RECT 0.498 0.213 0.526 0.215 ;
        RECT 0.146 0.638 0.535 0.666 ;
  END
END OAI21_X2_12T

MACRO OAI22_X1_12T
  CLASS core ;
  FOREIGN OAI22_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.672 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.199 0.27 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.279 0.398 0.576 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.192 0.206 0.512 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.192 0.08 0.576 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1409 0.638 0.306 0.666 ;
        RECT 0.306 0.182 0.334 0.638 ;
        RECT 0.306 0.638 0.334 0.666 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.101 0.37 0.131 ;
        RECT 0.37 0.101 0.398 0.131 ;
        RECT 0.37 0.131 0.398 0.211 ;
      LAYER M1 ;
        RECT 0.05 0.101 0.37 0.131 ;
        RECT 0.37 0.101 0.398 0.131 ;
        RECT 0.37 0.131 0.398 0.211 ;
  END
END OAI22_X1_12T

MACRO OAI22_X2_12T
  CLASS core ;
  FOREIGN OAI22_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.152 BY 1.152 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.256 0.462 0.279 ;
        RECT 0.434 0.279 0.462 0.466 ;
        RECT 0.434 0.466 0.462 0.494 ;
        RECT 0.462 0.466 0.6899 0.494 ;
        RECT 0.6899 0.279 0.718 0.466 ;
        RECT 0.6899 0.466 0.718 0.494 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.256 0.59 0.398 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.242 0.334 0.486 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.1419 0.512 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.386 0.27 0.53 ;
        RECT 0.242 0.53 0.27 0.558 ;
        RECT 0.27 0.53 0.37 0.558 ;
        RECT 0.37 0.169 0.398 0.197 ;
        RECT 0.37 0.197 0.398 0.278 ;
        RECT 0.37 0.278 0.398 0.386 ;
        RECT 0.37 0.386 0.398 0.53 ;
        RECT 0.37 0.53 0.398 0.558 ;
        RECT 0.398 0.169 0.626 0.197 ;
        RECT 0.398 0.53 0.626 0.558 ;
        RECT 0.626 0.169 0.654 0.197 ;
        RECT 0.626 0.197 0.654 0.278 ;
        RECT 0.626 0.53 0.654 0.558 ;
        RECT 0.654 0.53 0.6899 0.558 ;
        RECT 0.6899 0.53 0.718 0.558 ;
        RECT 0.6899 0.558 0.718 0.672 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.362 0.796 ;
        RECT 0.362 0.74 0.654 0.796 ;
        RECT 0.654 0.74 0.718 0.796 ;
        RECT 0.718 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.402 0.604 0.626 0.636 ;
        RECT 0.626 0.604 0.654 0.636 ;
        RECT 0.626 0.636 0.654 0.6959 ;
        RECT 0.041 0.099 0.6899 0.133 ;
        RECT 0.6899 0.099 0.718 0.133 ;
        RECT 0.6899 0.133 0.718 0.211 ;
        RECT 0.05 0.612 0.362 0.67 ;
      LAYER M1 ;
        RECT 0.402 0.604 0.626 0.636 ;
        RECT 0.626 0.604 0.654 0.636 ;
        RECT 0.626 0.636 0.654 0.6959 ;
        RECT 0.041 0.099 0.6899 0.133 ;
        RECT 0.6899 0.099 0.718 0.133 ;
        RECT 0.6899 0.133 0.718 0.211 ;
        RECT 0.05 0.612 0.362 0.67 ;
  END
END OAI22_X2_12T

MACRO OR2_X1_12T
  CLASS core ;
  FOREIGN OR2_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.096 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.243 0.078 0.641 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.114 0.334 0.64 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.13 0.1419 0.336 ;
        RECT 0.114 0.336 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.556 0.242 0.584 ;
        RECT 0.242 0.336 0.27 0.556 ;
        RECT 0.242 0.556 0.27 0.584 ;
      LAYER M1 ;
        RECT 0.114 0.13 0.1419 0.336 ;
        RECT 0.114 0.336 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.556 0.242 0.584 ;
        RECT 0.242 0.336 0.27 0.556 ;
        RECT 0.242 0.556 0.27 0.584 ;
  END
END OR2_X1_12T

MACRO OR2_X2_12T
  CLASS core ;
  FOREIGN OR2_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.672 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.1419 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.064 0.306 0.135 ;
        RECT 0.302 0.638 0.306 0.704 ;
        RECT 0.306 0.064 0.334 0.135 ;
        RECT 0.306 0.135 0.334 0.638 ;
        RECT 0.306 0.638 0.334 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.077 0.154 0.146 0.188 ;
        RECT 0.146 0.154 0.242 0.188 ;
        RECT 0.146 0.58 0.242 0.608 ;
        RECT 0.242 0.154 0.27 0.188 ;
        RECT 0.242 0.188 0.27 0.58 ;
        RECT 0.242 0.58 0.27 0.608 ;
      LAYER M1 ;
        RECT 0.077 0.154 0.146 0.188 ;
        RECT 0.146 0.154 0.242 0.188 ;
        RECT 0.146 0.58 0.242 0.608 ;
        RECT 0.242 0.154 0.27 0.188 ;
        RECT 0.242 0.188 0.27 0.58 ;
        RECT 0.242 0.58 0.27 0.608 ;
  END
END OR2_X2_12T

MACRO OR3_X1_12T
  CLASS core ;
  FOREIGN OR3_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.176 0.192 0.208 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.192 0.083 0.576 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.114 0.462 0.654 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.234 0.796 ;
        RECT 0.234 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.109 0.278 0.137 ;
        RECT 0.278 0.109 0.37 0.137 ;
        RECT 0.278 0.631 0.37 0.673 ;
        RECT 0.37 0.109 0.398 0.137 ;
        RECT 0.37 0.137 0.398 0.631 ;
        RECT 0.37 0.631 0.398 0.673 ;
        RECT 0.0859 0.636 0.234 0.668 ;
      LAYER M1 ;
        RECT 0.054 0.109 0.278 0.137 ;
        RECT 0.278 0.109 0.37 0.137 ;
        RECT 0.278 0.631 0.37 0.673 ;
        RECT 0.37 0.109 0.398 0.137 ;
        RECT 0.37 0.137 0.398 0.631 ;
        RECT 0.37 0.631 0.398 0.673 ;
        RECT 0.0859 0.636 0.234 0.668 ;
  END
END OR3_X1_12T

MACRO OR3_X2_12T
  CLASS core ;
  FOREIGN OR3_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.255 0.1419 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.526 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.231 0.27 0.448 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.366 0.064 0.37 0.13 ;
        RECT 0.366 0.636 0.37 0.704 ;
        RECT 0.37 0.064 0.398 0.13 ;
        RECT 0.37 0.13 0.398 0.636 ;
        RECT 0.37 0.636 0.398 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.302 0.796 ;
        RECT 0.302 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.5729 0.078 0.603 ;
        RECT 0.05 0.603 0.078 0.686 ;
        RECT 0.078 0.5729 0.302 0.603 ;
        RECT 0.06 0.155 0.1409 0.187 ;
        RECT 0.1409 0.155 0.306 0.187 ;
        RECT 0.1409 0.505 0.306 0.537 ;
        RECT 0.306 0.155 0.334 0.187 ;
        RECT 0.306 0.187 0.334 0.505 ;
        RECT 0.306 0.505 0.334 0.537 ;
      LAYER M1 ;
        RECT 0.05 0.5729 0.078 0.603 ;
        RECT 0.05 0.603 0.078 0.686 ;
        RECT 0.078 0.5729 0.302 0.603 ;
        RECT 0.06 0.155 0.1409 0.187 ;
        RECT 0.1409 0.155 0.306 0.187 ;
        RECT 0.1409 0.505 0.306 0.537 ;
        RECT 0.306 0.155 0.334 0.187 ;
        RECT 0.306 0.187 0.334 0.505 ;
        RECT 0.306 0.505 0.334 0.537 ;
  END
END OR3_X2_12T

MACRO OR4_X1_12T
  CLASS core ;
  FOREIGN OR4_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.192 0.272 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.198 0.1419 0.576 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.114 0.526 0.64 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.298 0.796 ;
        RECT 0.298 0.74 0.462 0.796 ;
        RECT 0.462 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.1019 0.338 0.13 ;
        RECT 0.338 0.1019 0.434 0.13 ;
        RECT 0.338 0.63 0.434 0.662 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.63 ;
        RECT 0.434 0.63 0.462 0.662 ;
        RECT 0.146 0.617 0.298 0.655 ;
      LAYER M1 ;
        RECT 0.054 0.1019 0.338 0.13 ;
        RECT 0.338 0.1019 0.434 0.13 ;
        RECT 0.338 0.63 0.434 0.662 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.63 ;
        RECT 0.434 0.63 0.462 0.662 ;
        RECT 0.146 0.617 0.298 0.655 ;
  END
END OR4_X1_12T

MACRO OR4_X2_12T
  CLASS core ;
  FOREIGN OR4_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.96 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.53 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.213 0.27 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.213 0.1419 0.576 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.191 0.078 0.576 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.496 0.128 0.528 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.302 0.796 ;
        RECT 0.302 0.74 0.46 0.796 ;
        RECT 0.46 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.146 0.623 0.302 0.681 ;
        RECT 0.054 0.0869 0.342 0.145 ;
        RECT 0.342 0.0869 0.432 0.145 ;
        RECT 0.342 0.5679 0.432 0.624 ;
        RECT 0.432 0.0869 0.46 0.145 ;
        RECT 0.432 0.145 0.46 0.5679 ;
        RECT 0.432 0.5679 0.46 0.624 ;
      LAYER M1 ;
        RECT 0.146 0.623 0.302 0.681 ;
        RECT 0.054 0.0869 0.342 0.145 ;
        RECT 0.342 0.0869 0.432 0.145 ;
        RECT 0.342 0.5679 0.432 0.624 ;
        RECT 0.432 0.0869 0.46 0.145 ;
        RECT 0.432 0.145 0.46 0.5679 ;
        RECT 0.432 0.5679 0.46 0.624 ;
  END
END OR4_X2_12T

MACRO SDFFRNQ_X1_12T
  CLASS core ;
  FOREIGN SDFFRNQ_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.88 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.363 0.515 0.528 ;
        RECT 0.515 0.363 0.526 0.528 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.965 0.338 1.454 0.366 ;
        RECT 1.454 0.338 1.592 0.366 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.372 0.334 0.5719 ;
        RECT 0.306 0.5719 0.334 0.6 ;
        RECT 0.334 0.5719 0.515 0.6 ;
        RECT 0.515 0.5719 0.562 0.6 ;
        RECT 0.562 0.314 0.59 0.372 ;
        RECT 0.562 0.372 0.59 0.5719 ;
        RECT 0.562 0.5719 0.59 0.6 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.363 0.398 0.512 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.276 0.078 0.534 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.064 1.872 0.704 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.754 0.796 ;
        RECT 0.754 0.74 0.782 0.796 ;
        RECT 0.782 0.74 1.066 0.796 ;
        RECT 1.066 0.74 1.422 0.796 ;
        RECT 1.422 0.74 1.49 0.796 ;
        RECT 1.49 0.74 1.742 0.796 ;
        RECT 1.742 0.74 1.93 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.93 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.53 1.326 0.558 ;
        RECT 0.722 0.402 1.121 0.43 ;
        RECT 0.082 0.274 1.454 0.302 ;
      LAYER MINT1 ;
        RECT 0.146 0.53 1.326 0.558 ;
        RECT 0.722 0.402 1.121 0.43 ;
        RECT 0.082 0.274 1.454 0.302 ;
      LAYER M1 ;
        RECT 0.045 0.096 0.083 0.2039 ;
        RECT 0.045 0.2039 0.083 0.232 ;
        RECT 0.045 0.604 0.083 0.632 ;
        RECT 0.045 0.632 0.083 0.6879 ;
        RECT 0.083 0.2039 0.114 0.232 ;
        RECT 0.083 0.604 0.114 0.632 ;
        RECT 0.114 0.2039 0.1419 0.232 ;
        RECT 0.114 0.232 0.1419 0.604 ;
        RECT 0.114 0.604 0.1419 0.632 ;
        RECT 0.242 0.096 0.27 0.267 ;
        RECT 0.242 0.267 0.27 0.295 ;
        RECT 0.242 0.295 0.27 0.672 ;
        RECT 0.27 0.267 0.515 0.295 ;
        RECT 0.338 0.184 0.626 0.212 ;
        RECT 0.626 0.184 0.654 0.212 ;
        RECT 0.626 0.212 0.654 0.276 ;
        RECT 0.392 0.636 0.754 0.668 ;
        RECT 0.754 0.247 0.782 0.546 ;
        RECT 0.466 0.1019 0.878 0.13 ;
        RECT 1.061 0.24 1.098 0.446 ;
        RECT 1.202 0.171 1.23 0.511 ;
        RECT 1.458 0.146 1.49 0.6979 ;
        RECT 1.165 0.618 1.33 0.646 ;
        RECT 1.33 0.064 1.358 0.092 ;
        RECT 1.33 0.092 1.358 0.366 ;
        RECT 1.33 0.366 1.358 0.618 ;
        RECT 1.33 0.618 1.358 0.646 ;
        RECT 1.358 0.064 1.607 0.092 ;
        RECT 1.607 0.064 1.635 0.092 ;
        RECT 1.607 0.092 1.635 0.366 ;
        RECT 1.554 0.46 1.582 0.624 ;
        RECT 1.554 0.624 1.582 0.68 ;
        RECT 1.582 0.624 1.714 0.68 ;
        RECT 1.714 0.072 1.742 0.46 ;
        RECT 1.714 0.46 1.742 0.624 ;
        RECT 1.714 0.624 1.742 0.68 ;
        RECT 0.178 0.125 0.206 0.574 ;
        RECT 0.6899 0.387 0.718 0.59 ;
        RECT 0.8179 0.257 0.85 0.469 ;
        RECT 0.6899 0.166 0.718 0.194 ;
        RECT 0.6899 0.194 0.718 0.276 ;
        RECT 0.718 0.166 0.942 0.194 ;
        RECT 0.991 0.242 1.025 0.422 ;
        RECT 0.79 0.636 1.066 0.668 ;
        RECT 0.904 0.274 0.932 0.49 ;
        RECT 0.904 0.49 0.932 0.518 ;
        RECT 0.932 0.49 1.1339 0.518 ;
        RECT 1.1339 0.082 1.166 0.274 ;
        RECT 1.1339 0.274 1.166 0.49 ;
        RECT 1.1339 0.49 1.166 0.518 ;
        RECT 1.266 0.178 1.294 0.574 ;
        RECT 1.3939 0.178 1.422 0.494 ;
        RECT 1.532 0.154 1.571 0.416 ;
      LAYER V1 ;
        RECT 0.114 0.274 0.1419 0.302 ;
        RECT 0.178 0.53 0.206 0.558 ;
        RECT 0.6899 0.53 0.718 0.558 ;
        RECT 0.754 0.402 0.782 0.43 ;
        RECT 0.8179 0.274 0.846 0.302 ;
        RECT 0.997 0.338 1.025 0.366 ;
        RECT 1.061 0.402 1.089 0.43 ;
        RECT 1.202 0.274 1.23 0.302 ;
        RECT 1.266 0.53 1.294 0.558 ;
        RECT 1.3939 0.274 1.422 0.302 ;
        RECT 1.532 0.338 1.56 0.366 ;
      LAYER M1 ;
        RECT 0.045 0.096 0.083 0.2039 ;
        RECT 0.045 0.2039 0.083 0.232 ;
        RECT 0.045 0.604 0.083 0.632 ;
        RECT 0.045 0.632 0.083 0.6879 ;
        RECT 0.083 0.2039 0.114 0.232 ;
        RECT 0.083 0.604 0.114 0.632 ;
        RECT 0.114 0.2039 0.1419 0.232 ;
        RECT 0.114 0.232 0.1419 0.604 ;
        RECT 0.114 0.604 0.1419 0.632 ;
        RECT 0.242 0.096 0.27 0.267 ;
        RECT 0.242 0.267 0.27 0.295 ;
        RECT 0.242 0.295 0.27 0.672 ;
        RECT 0.27 0.267 0.515 0.295 ;
        RECT 0.338 0.184 0.626 0.212 ;
        RECT 0.626 0.184 0.654 0.212 ;
        RECT 0.626 0.212 0.654 0.276 ;
        RECT 0.392 0.636 0.754 0.668 ;
        RECT 0.754 0.247 0.782 0.546 ;
        RECT 0.466 0.1019 0.878 0.13 ;
        RECT 1.061 0.24 1.098 0.446 ;
        RECT 1.202 0.171 1.23 0.511 ;
        RECT 1.458 0.146 1.49 0.6979 ;
        RECT 1.165 0.618 1.33 0.646 ;
        RECT 1.33 0.064 1.358 0.092 ;
        RECT 1.33 0.092 1.358 0.366 ;
        RECT 1.33 0.366 1.358 0.618 ;
        RECT 1.33 0.618 1.358 0.646 ;
        RECT 1.358 0.064 1.607 0.092 ;
        RECT 1.607 0.064 1.635 0.092 ;
        RECT 1.607 0.092 1.635 0.366 ;
        RECT 1.554 0.46 1.582 0.624 ;
        RECT 1.554 0.624 1.582 0.68 ;
        RECT 1.582 0.624 1.714 0.68 ;
        RECT 1.714 0.072 1.742 0.46 ;
        RECT 1.714 0.46 1.742 0.624 ;
        RECT 1.714 0.624 1.742 0.68 ;
        RECT 0.178 0.125 0.206 0.574 ;
        RECT 0.6899 0.387 0.718 0.59 ;
        RECT 0.8179 0.257 0.85 0.469 ;
        RECT 0.6899 0.166 0.718 0.194 ;
        RECT 0.6899 0.194 0.718 0.276 ;
        RECT 0.718 0.166 0.942 0.194 ;
        RECT 0.991 0.242 1.025 0.422 ;
        RECT 0.79 0.636 1.066 0.668 ;
        RECT 0.904 0.274 0.932 0.49 ;
        RECT 0.904 0.49 0.932 0.518 ;
        RECT 0.932 0.49 1.1339 0.518 ;
        RECT 1.1339 0.082 1.166 0.274 ;
        RECT 1.1339 0.274 1.166 0.49 ;
        RECT 1.1339 0.49 1.166 0.518 ;
        RECT 1.266 0.178 1.294 0.574 ;
        RECT 1.3939 0.178 1.422 0.494 ;
        RECT 1.532 0.154 1.571 0.416 ;
  END
END SDFFRNQ_X1_12T

MACRO SDFFSNQ_X1_12T
  CLASS core ;
  FOREIGN SDFFSNQ_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.88 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.384 0.51 0.528 ;
        RECT 0.51 0.384 0.526 0.528 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.372 0.334 0.5719 ;
        RECT 0.306 0.5719 0.334 0.6 ;
        RECT 0.334 0.5719 0.51 0.6 ;
        RECT 0.51 0.5719 0.562 0.6 ;
        RECT 0.562 0.314 0.59 0.372 ;
        RECT 0.562 0.372 0.59 0.5719 ;
        RECT 0.562 0.5719 0.59 0.6 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.363 0.398 0.512 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.958 0.338 1.454 0.366 ;
        RECT 1.454 0.338 1.586 0.366 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.272 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.064 1.872 0.704 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.746 0.796 ;
        RECT 0.746 0.74 0.782 0.796 ;
        RECT 0.782 0.74 0.862 0.796 ;
        RECT 0.862 0.74 1.646 0.796 ;
        RECT 1.646 0.74 1.742 0.796 ;
        RECT 1.742 0.74 1.93 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.93 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.53 1.326 0.558 ;
        RECT 0.722 0.402 1.114 0.43 ;
        RECT 0.082 0.274 1.454 0.302 ;
      LAYER MINT1 ;
        RECT 0.146 0.53 1.326 0.558 ;
        RECT 0.722 0.402 1.114 0.43 ;
        RECT 0.082 0.274 1.454 0.302 ;
      LAYER M1 ;
        RECT 0.048 0.064 0.08 0.2 ;
        RECT 0.048 0.2 0.08 0.228 ;
        RECT 0.048 0.604 0.08 0.632 ;
        RECT 0.048 0.632 0.08 0.6879 ;
        RECT 0.08 0.2 0.114 0.228 ;
        RECT 0.08 0.604 0.114 0.632 ;
        RECT 0.114 0.2 0.1419 0.228 ;
        RECT 0.114 0.228 0.1419 0.604 ;
        RECT 0.114 0.604 0.1419 0.632 ;
        RECT 0.242 0.082 0.27 0.266 ;
        RECT 0.242 0.266 0.27 0.295 ;
        RECT 0.242 0.295 0.27 0.296 ;
        RECT 0.242 0.296 0.27 0.686 ;
        RECT 0.27 0.266 0.434 0.295 ;
        RECT 0.434 0.266 0.51 0.295 ;
        RECT 0.434 0.295 0.51 0.296 ;
        RECT 0.338 0.184 0.626 0.212 ;
        RECT 0.626 0.184 0.654 0.212 ;
        RECT 0.626 0.212 0.654 0.276 ;
        RECT 0.392 0.636 0.746 0.668 ;
        RECT 0.754 0.238 0.782 0.547 ;
        RECT 0.466 0.1019 0.878 0.13 ;
        RECT 0.98 0.322 1.018 0.419 ;
        RECT 0.898 0.274 0.926 0.487 ;
        RECT 0.898 0.487 0.926 0.515 ;
        RECT 0.926 0.487 1.008 0.515 ;
        RECT 1.008 0.487 1.04 0.515 ;
        RECT 1.008 0.515 1.04 0.704 ;
        RECT 1.04 0.487 1.1379 0.515 ;
        RECT 1.1379 0.098 1.166 0.274 ;
        RECT 1.1379 0.274 1.166 0.487 ;
        RECT 1.1379 0.487 1.166 0.515 ;
        RECT 1.266 0.178 1.294 0.574 ;
        RECT 1.3939 0.178 1.422 0.402 ;
        RECT 1.526 0.184 1.554 0.403 ;
        RECT 1.402 0.638 1.646 0.666 ;
        RECT 0.178 0.096 0.206 0.619 ;
        RECT 0.654 0.387 0.682 0.574 ;
        RECT 0.83 0.257 0.862 0.469 ;
        RECT 0.6899 0.166 0.718 0.194 ;
        RECT 0.6899 0.194 0.718 0.276 ;
        RECT 0.718 0.166 0.942 0.194 ;
        RECT 1.054 0.24 1.092 0.446 ;
        RECT 1.202 0.171 1.23 0.383 ;
        RECT 1.165 0.618 1.33 0.646 ;
        RECT 1.33 0.082 1.358 0.11 ;
        RECT 1.33 0.11 1.358 0.366 ;
        RECT 1.33 0.366 1.358 0.618 ;
        RECT 1.33 0.618 1.358 0.646 ;
        RECT 1.358 0.082 1.607 0.11 ;
        RECT 1.607 0.082 1.645 0.11 ;
        RECT 1.607 0.11 1.645 0.366 ;
        RECT 1.462 0.402 1.49 0.574 ;
        RECT 1.462 0.574 1.49 0.602 ;
        RECT 1.49 0.574 1.714 0.602 ;
        RECT 1.714 0.096 1.742 0.402 ;
        RECT 1.714 0.402 1.742 0.574 ;
        RECT 1.714 0.574 1.742 0.602 ;
      LAYER V1 ;
        RECT 0.114 0.274 0.1419 0.302 ;
        RECT 0.178 0.53 0.206 0.558 ;
        RECT 0.654 0.53 0.682 0.558 ;
        RECT 0.754 0.402 0.782 0.43 ;
        RECT 0.834 0.274 0.862 0.302 ;
        RECT 0.99 0.338 1.018 0.366 ;
        RECT 1.054 0.402 1.082 0.43 ;
        RECT 1.202 0.274 1.23 0.302 ;
        RECT 1.266 0.53 1.294 0.558 ;
        RECT 1.3939 0.274 1.422 0.302 ;
        RECT 1.526 0.338 1.554 0.366 ;
      LAYER M1 ;
        RECT 0.048 0.064 0.08 0.2 ;
        RECT 0.048 0.2 0.08 0.228 ;
        RECT 0.048 0.604 0.08 0.632 ;
        RECT 0.048 0.632 0.08 0.6879 ;
        RECT 0.08 0.2 0.114 0.228 ;
        RECT 0.08 0.604 0.114 0.632 ;
        RECT 0.114 0.2 0.1419 0.228 ;
        RECT 0.114 0.228 0.1419 0.604 ;
        RECT 0.114 0.604 0.1419 0.632 ;
        RECT 0.242 0.082 0.27 0.266 ;
        RECT 0.242 0.266 0.27 0.295 ;
        RECT 0.242 0.295 0.27 0.296 ;
        RECT 0.242 0.296 0.27 0.686 ;
        RECT 0.27 0.266 0.434 0.295 ;
        RECT 0.434 0.266 0.51 0.295 ;
        RECT 0.434 0.295 0.51 0.296 ;
        RECT 0.338 0.184 0.626 0.212 ;
        RECT 0.626 0.184 0.654 0.212 ;
        RECT 0.626 0.212 0.654 0.276 ;
        RECT 0.392 0.636 0.746 0.668 ;
        RECT 0.754 0.238 0.782 0.547 ;
        RECT 0.466 0.1019 0.878 0.13 ;
        RECT 0.98 0.322 1.018 0.419 ;
        RECT 0.898 0.274 0.926 0.487 ;
        RECT 0.898 0.487 0.926 0.515 ;
        RECT 0.926 0.487 1.008 0.515 ;
        RECT 1.008 0.487 1.04 0.515 ;
        RECT 1.008 0.515 1.04 0.704 ;
        RECT 1.04 0.487 1.1379 0.515 ;
        RECT 1.1379 0.098 1.166 0.274 ;
        RECT 1.1379 0.274 1.166 0.487 ;
        RECT 1.1379 0.487 1.166 0.515 ;
        RECT 1.266 0.178 1.294 0.574 ;
        RECT 1.3939 0.178 1.422 0.402 ;
        RECT 1.526 0.184 1.554 0.403 ;
        RECT 1.402 0.638 1.646 0.666 ;
        RECT 0.178 0.096 0.206 0.619 ;
        RECT 0.654 0.387 0.682 0.574 ;
        RECT 0.83 0.257 0.862 0.469 ;
        RECT 0.6899 0.166 0.718 0.194 ;
        RECT 0.6899 0.194 0.718 0.276 ;
        RECT 0.718 0.166 0.942 0.194 ;
        RECT 1.054 0.24 1.092 0.446 ;
        RECT 1.202 0.171 1.23 0.383 ;
        RECT 1.165 0.618 1.33 0.646 ;
        RECT 1.33 0.082 1.358 0.11 ;
        RECT 1.33 0.11 1.358 0.366 ;
        RECT 1.33 0.366 1.358 0.618 ;
        RECT 1.33 0.618 1.358 0.646 ;
        RECT 1.358 0.082 1.607 0.11 ;
        RECT 1.607 0.082 1.645 0.11 ;
        RECT 1.607 0.11 1.645 0.366 ;
        RECT 1.462 0.402 1.49 0.574 ;
        RECT 1.462 0.574 1.49 0.602 ;
        RECT 1.49 0.574 1.714 0.602 ;
        RECT 1.714 0.096 1.742 0.402 ;
        RECT 1.714 0.402 1.742 0.574 ;
        RECT 1.714 0.574 1.742 0.602 ;
  END
END SDFFSNQ_X1_12T

MACRO TBUF_X1_12T
  CLASS core ;
  FOREIGN TBUF_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.056 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.492 ;
        RECT 0.114 0.492 0.1419 0.52 ;
        RECT 0.1419 0.492 0.206 0.52 ;
        RECT 0.206 0.492 0.242 0.52 ;
        RECT 0.242 0.306 0.27 0.384 ;
        RECT 0.242 0.384 0.27 0.492 ;
        RECT 0.242 0.492 0.27 0.52 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.37 0.462 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.064 0.656 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.588 0.796 ;
        RECT 0.588 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.418 ;
        RECT 0.05 0.418 0.078 0.686 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.418 ;
        RECT 0.146 0.574 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.574 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.574 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.314 ;
        RECT 0.306 0.314 0.334 0.574 ;
        RECT 0.306 0.574 0.334 0.602 ;
        RECT 0.334 0.1019 0.51 0.13 ;
        RECT 0.51 0.1019 0.542 0.13 ;
        RECT 0.51 0.13 0.542 0.23 ;
        RECT 0.51 0.23 0.542 0.258 ;
        RECT 0.51 0.258 0.542 0.314 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.376 ;
        RECT 0.37 0.376 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.56 0.666 ;
        RECT 0.56 0.376 0.588 0.638 ;
        RECT 0.56 0.638 0.588 0.666 ;
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.418 ;
        RECT 0.05 0.418 0.078 0.686 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.418 ;
        RECT 0.146 0.574 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.574 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.574 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.314 ;
        RECT 0.306 0.314 0.334 0.574 ;
        RECT 0.306 0.574 0.334 0.602 ;
        RECT 0.334 0.1019 0.51 0.13 ;
        RECT 0.51 0.1019 0.542 0.13 ;
        RECT 0.51 0.13 0.542 0.23 ;
        RECT 0.51 0.23 0.542 0.258 ;
        RECT 0.51 0.258 0.542 0.314 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.376 ;
        RECT 0.37 0.376 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.56 0.666 ;
        RECT 0.56 0.376 0.588 0.638 ;
        RECT 0.56 0.638 0.588 0.666 ;
  END
END TBUF_X1_12T

MACRO TBUF_X2_12T
  CLASS core ;
  FOREIGN TBUF_X2_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.152 BY 1.152 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.504 ;
        RECT 0.114 0.504 0.1419 0.532 ;
        RECT 0.1419 0.504 0.206 0.532 ;
        RECT 0.206 0.504 0.242 0.532 ;
        RECT 0.242 0.306 0.27 0.384 ;
        RECT 0.242 0.384 0.27 0.504 ;
        RECT 0.242 0.504 0.27 0.532 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.382 0.462 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.07 0.656 0.6959 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.53 0.796 ;
        RECT 0.53 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.612 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.146 0.5679 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.5679 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.5679 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.314 ;
        RECT 0.306 0.314 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.602 ;
        RECT 0.334 0.1019 0.482 0.13 ;
        RECT 0.482 0.1019 0.514 0.13 ;
        RECT 0.482 0.13 0.514 0.23 ;
        RECT 0.482 0.23 0.514 0.258 ;
        RECT 0.482 0.258 0.514 0.314 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.443 ;
        RECT 0.37 0.443 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.498 0.666 ;
        RECT 0.498 0.443 0.53 0.638 ;
        RECT 0.498 0.638 0.53 0.666 ;
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.612 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.146 0.5679 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.5679 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.5679 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.314 ;
        RECT 0.306 0.314 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.602 ;
        RECT 0.334 0.1019 0.482 0.13 ;
        RECT 0.482 0.1019 0.514 0.13 ;
        RECT 0.482 0.13 0.514 0.23 ;
        RECT 0.482 0.23 0.514 0.258 ;
        RECT 0.482 0.258 0.514 0.314 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.443 ;
        RECT 0.37 0.443 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.498 0.666 ;
        RECT 0.498 0.443 0.53 0.638 ;
        RECT 0.498 0.638 0.53 0.666 ;
  END
END TBUF_X2_12T

MACRO TBUF_X4_12T
  CLASS core ;
  FOREIGN TBUF_X4_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.44 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.484 ;
        RECT 0.114 0.484 0.1419 0.512 ;
        RECT 0.1419 0.484 0.206 0.512 ;
        RECT 0.206 0.484 0.242 0.512 ;
        RECT 0.242 0.306 0.27 0.384 ;
        RECT 0.242 0.384 0.27 0.484 ;
        RECT 0.242 0.484 0.27 0.512 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.3459 0.462 0.594 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.6879 0.064 0.72 0.224 ;
        RECT 0.6879 0.224 0.72 0.256 ;
        RECT 0.6879 0.512 0.72 0.54 ;
        RECT 0.6879 0.54 0.72 0.5709 ;
        RECT 0.6879 0.5709 0.72 0.704 ;
        RECT 0.72 0.224 0.8129 0.256 ;
        RECT 0.72 0.512 0.8129 0.54 ;
        RECT 0.8129 0.064 0.8139 0.224 ;
        RECT 0.8129 0.224 0.8139 0.256 ;
        RECT 0.8129 0.512 0.8139 0.54 ;
        RECT 0.8139 0.064 0.8159 0.224 ;
        RECT 0.8139 0.224 0.8159 0.256 ;
        RECT 0.8139 0.512 0.8159 0.54 ;
        RECT 0.8159 0.064 0.838 0.224 ;
        RECT 0.8159 0.224 0.838 0.256 ;
        RECT 0.8159 0.512 0.838 0.54 ;
        RECT 0.8159 0.54 0.838 0.5709 ;
        RECT 0.8159 0.5709 0.838 0.704 ;
        RECT 0.838 0.064 0.848 0.224 ;
        RECT 0.838 0.224 0.848 0.256 ;
        RECT 0.838 0.512 0.848 0.54 ;
        RECT 0.838 0.54 0.848 0.5709 ;
        RECT 0.838 0.5709 0.848 0.704 ;
        RECT 0.848 0.064 0.851 0.224 ;
        RECT 0.848 0.224 0.851 0.256 ;
        RECT 0.848 0.512 0.851 0.54 ;
        RECT 0.848 0.54 0.851 0.5709 ;
        RECT 0.851 0.224 0.882 0.256 ;
        RECT 0.851 0.512 0.882 0.54 ;
        RECT 0.851 0.54 0.882 0.5709 ;
        RECT 0.882 0.224 0.91 0.256 ;
        RECT 0.882 0.256 0.91 0.512 ;
        RECT 0.882 0.512 0.91 0.54 ;
        RECT 0.882 0.54 0.91 0.5709 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.8139 0.796 ;
        RECT 0.8139 0.74 0.838 0.796 ;
        RECT 0.838 0.74 0.97 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.97 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.388 ;
        RECT 0.37 0.388 0.398 0.414 ;
        RECT 0.37 0.414 0.398 0.458 ;
        RECT 0.37 0.458 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.526 0.666 ;
        RECT 0.526 0.388 0.582 0.414 ;
        RECT 0.526 0.414 0.582 0.458 ;
        RECT 0.526 0.458 0.582 0.638 ;
        RECT 0.526 0.638 0.582 0.666 ;
        RECT 0.582 0.414 0.8139 0.458 ;
        RECT 0.05 0.096 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.594 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.146 0.5679 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.5679 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.5679 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.292 ;
        RECT 0.306 0.292 0.334 0.32 ;
        RECT 0.306 0.32 0.334 0.352 ;
        RECT 0.306 0.352 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.602 ;
        RECT 0.334 0.1019 0.526 0.13 ;
        RECT 0.526 0.1019 0.582 0.13 ;
        RECT 0.526 0.13 0.582 0.23 ;
        RECT 0.526 0.23 0.582 0.258 ;
        RECT 0.526 0.258 0.582 0.292 ;
        RECT 0.526 0.292 0.582 0.32 ;
        RECT 0.526 0.32 0.582 0.352 ;
        RECT 0.582 0.292 0.838 0.32 ;
      LAYER M1 ;
        RECT 0.082 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.388 ;
        RECT 0.37 0.388 0.398 0.414 ;
        RECT 0.37 0.414 0.398 0.458 ;
        RECT 0.37 0.458 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.526 0.666 ;
        RECT 0.526 0.388 0.582 0.414 ;
        RECT 0.526 0.414 0.582 0.458 ;
        RECT 0.526 0.458 0.582 0.638 ;
        RECT 0.526 0.638 0.582 0.666 ;
        RECT 0.582 0.414 0.8139 0.458 ;
        RECT 0.05 0.096 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.594 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.146 0.5679 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.5679 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.5679 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.292 ;
        RECT 0.306 0.292 0.334 0.32 ;
        RECT 0.306 0.32 0.334 0.352 ;
        RECT 0.306 0.352 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.602 ;
        RECT 0.334 0.1019 0.526 0.13 ;
        RECT 0.526 0.1019 0.582 0.13 ;
        RECT 0.526 0.13 0.582 0.23 ;
        RECT 0.526 0.23 0.582 0.258 ;
        RECT 0.526 0.258 0.582 0.292 ;
        RECT 0.526 0.292 0.582 0.32 ;
        RECT 0.526 0.32 0.582 0.352 ;
        RECT 0.582 0.292 0.838 0.32 ;
  END
END TBUF_X4_12T

MACRO TBUF_X8_12T
  CLASS core ;
  FOREIGN TBUF_X8_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.016 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.484 ;
        RECT 0.114 0.484 0.1419 0.512 ;
        RECT 0.1419 0.484 0.222 0.512 ;
        RECT 0.222 0.484 0.306 0.512 ;
        RECT 0.306 0.32 0.334 0.384 ;
        RECT 0.306 0.384 0.334 0.484 ;
        RECT 0.306 0.484 0.334 0.512 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.3459 0.526 0.402 ;
        RECT 0.498 0.402 0.526 0.434 ;
        RECT 0.498 0.434 0.526 0.576 ;
        RECT 0.526 0.402 0.622 0.434 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8159 0.064 0.848 0.133 ;
        RECT 0.8159 0.133 0.848 0.16 ;
        RECT 0.8159 0.16 0.848 0.192 ;
        RECT 0.8159 0.519 0.848 0.577 ;
        RECT 0.8159 0.577 0.848 0.578 ;
        RECT 0.8159 0.578 0.848 0.704 ;
        RECT 0.848 0.16 1.183 0.192 ;
        RECT 0.848 0.519 1.183 0.577 ;
        RECT 1.183 0.16 1.198 0.192 ;
        RECT 1.183 0.519 1.198 0.577 ;
        RECT 1.198 0.16 1.2 0.192 ;
        RECT 1.198 0.519 1.2 0.577 ;
        RECT 1.2 0.064 1.232 0.133 ;
        RECT 1.2 0.133 1.232 0.16 ;
        RECT 1.2 0.16 1.232 0.192 ;
        RECT 1.2 0.519 1.232 0.577 ;
        RECT 1.2 0.577 1.232 0.578 ;
        RECT 1.2 0.578 1.232 0.704 ;
        RECT 1.232 0.133 1.266 0.16 ;
        RECT 1.232 0.16 1.266 0.192 ;
        RECT 1.232 0.519 1.266 0.577 ;
        RECT 1.232 0.577 1.266 0.578 ;
        RECT 1.266 0.133 1.294 0.16 ;
        RECT 1.266 0.16 1.294 0.192 ;
        RECT 1.266 0.192 1.294 0.519 ;
        RECT 1.266 0.519 1.294 0.577 ;
        RECT 1.266 0.577 1.294 0.578 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.183 0.796 ;
        RECT 1.183 0.74 1.198 0.796 ;
        RECT 1.198 0.74 1.354 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.354 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.43 ;
        RECT 0.05 0.43 0.078 0.638 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.222 0.34 ;
        RECT 0.178 0.34 0.222 0.43 ;
        RECT 0.146 0.574 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.574 0.23 0.602 ;
        RECT 0.23 0.1019 0.37 0.13 ;
        RECT 0.23 0.23 0.37 0.258 ;
        RECT 0.23 0.574 0.37 0.602 ;
        RECT 0.37 0.1019 0.398 0.13 ;
        RECT 0.37 0.23 0.398 0.258 ;
        RECT 0.37 0.258 0.398 0.2859 ;
        RECT 0.37 0.2859 0.398 0.342 ;
        RECT 0.37 0.342 0.398 0.574 ;
        RECT 0.37 0.574 0.398 0.602 ;
        RECT 0.398 0.1019 0.6899 0.13 ;
        RECT 0.6899 0.1019 0.718 0.13 ;
        RECT 0.6899 0.13 0.718 0.23 ;
        RECT 0.6899 0.23 0.718 0.258 ;
        RECT 0.6899 0.258 0.718 0.2859 ;
        RECT 0.6899 0.2859 0.718 0.342 ;
        RECT 0.718 0.258 1.198 0.2859 ;
        RECT 0.122 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.434 0.194 ;
        RECT 0.274 0.638 0.434 0.666 ;
        RECT 0.434 0.166 0.462 0.194 ;
        RECT 0.434 0.194 0.462 0.386 ;
        RECT 0.434 0.386 0.462 0.403 ;
        RECT 0.434 0.403 0.462 0.461 ;
        RECT 0.434 0.461 0.462 0.638 ;
        RECT 0.434 0.638 0.462 0.666 ;
        RECT 0.462 0.638 0.66 0.666 ;
        RECT 0.66 0.386 0.718 0.403 ;
        RECT 0.66 0.403 0.718 0.461 ;
        RECT 0.66 0.461 0.718 0.638 ;
        RECT 0.66 0.638 0.718 0.666 ;
        RECT 0.718 0.403 1.183 0.461 ;
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.43 ;
        RECT 0.05 0.43 0.078 0.638 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.222 0.34 ;
        RECT 0.178 0.34 0.222 0.43 ;
        RECT 0.146 0.574 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.574 0.23 0.602 ;
        RECT 0.23 0.1019 0.37 0.13 ;
        RECT 0.23 0.23 0.37 0.258 ;
        RECT 0.23 0.574 0.37 0.602 ;
        RECT 0.37 0.1019 0.398 0.13 ;
        RECT 0.37 0.23 0.398 0.258 ;
        RECT 0.37 0.258 0.398 0.2859 ;
        RECT 0.37 0.2859 0.398 0.342 ;
        RECT 0.37 0.342 0.398 0.574 ;
        RECT 0.37 0.574 0.398 0.602 ;
        RECT 0.398 0.1019 0.6899 0.13 ;
        RECT 0.6899 0.1019 0.718 0.13 ;
        RECT 0.6899 0.13 0.718 0.23 ;
        RECT 0.6899 0.23 0.718 0.258 ;
        RECT 0.6899 0.258 0.718 0.2859 ;
        RECT 0.6899 0.2859 0.718 0.342 ;
        RECT 0.718 0.258 1.198 0.2859 ;
        RECT 0.122 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.434 0.194 ;
        RECT 0.274 0.638 0.434 0.666 ;
        RECT 0.434 0.166 0.462 0.194 ;
        RECT 0.434 0.194 0.462 0.386 ;
        RECT 0.434 0.386 0.462 0.403 ;
        RECT 0.434 0.403 0.462 0.461 ;
        RECT 0.434 0.461 0.462 0.638 ;
        RECT 0.434 0.638 0.462 0.666 ;
        RECT 0.462 0.638 0.66 0.666 ;
        RECT 0.66 0.386 0.718 0.403 ;
        RECT 0.66 0.403 0.718 0.461 ;
        RECT 0.66 0.461 0.718 0.638 ;
        RECT 0.66 0.638 0.718 0.666 ;
        RECT 0.718 0.403 1.183 0.461 ;
  END
END TBUF_X8_12T

MACRO TBUF_X12_12T
  CLASS core ;
  FOREIGN TBUF_X12_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.592 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.51 ;
        RECT 0.114 0.51 0.1419 0.538 ;
        RECT 0.1419 0.51 0.206 0.538 ;
        RECT 0.206 0.51 0.242 0.538 ;
        RECT 0.242 0.306 0.27 0.384 ;
        RECT 0.242 0.384 0.27 0.51 ;
        RECT 0.242 0.51 0.27 0.538 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.402 0.498 0.448 ;
        RECT 0.498 0.3459 0.526 0.402 ;
        RECT 0.498 0.402 0.526 0.448 ;
        RECT 0.526 0.402 0.626 0.448 ;
        RECT 0.626 0.402 0.654 0.448 ;
        RECT 0.626 0.448 0.654 0.576 ;
        RECT 0.654 0.402 0.71 0.448 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.684 0.796 ;
        RECT 1.684 0.74 1.738 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.738 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.356 ;
        RECT 0.37 0.356 0.398 0.378 ;
        RECT 0.37 0.378 0.398 0.426 ;
        RECT 0.37 0.426 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.783 0.666 ;
        RECT 0.783 0.356 0.839 0.378 ;
        RECT 0.783 0.378 0.839 0.426 ;
        RECT 0.783 0.426 0.839 0.638 ;
        RECT 0.783 0.638 0.839 0.666 ;
        RECT 0.839 0.378 1.557 0.426 ;
        RECT 0.882 0.1019 0.931 0.13 ;
        RECT 0.931 0.1019 0.989 0.13 ;
        RECT 0.931 0.532 0.989 0.5639 ;
        RECT 0.931 0.5639 0.989 0.62 ;
        RECT 0.989 0.1019 1.572 0.13 ;
        RECT 0.989 0.532 1.572 0.5639 ;
        RECT 1.572 0.073 1.586 0.1019 ;
        RECT 1.572 0.1019 1.586 0.13 ;
        RECT 1.572 0.532 1.586 0.5639 ;
        RECT 1.586 0.073 1.614 0.1019 ;
        RECT 1.586 0.1019 1.614 0.13 ;
        RECT 1.586 0.532 1.614 0.5639 ;
        RECT 1.586 0.5639 1.614 0.62 ;
        RECT 1.586 0.62 1.614 0.624 ;
        RECT 1.614 0.073 1.6279 0.1019 ;
        RECT 1.614 0.1019 1.6279 0.13 ;
        RECT 1.614 0.532 1.6279 0.5639 ;
        RECT 1.6279 0.1019 1.629 0.13 ;
        RECT 1.6279 0.532 1.629 0.5639 ;
        RECT 1.629 0.1019 1.684 0.13 ;
        RECT 1.629 0.13 1.684 0.532 ;
        RECT 1.629 0.532 1.684 0.5639 ;
        RECT 0.05 0.1739 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.672 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.1419 0.1019 0.146 0.13 ;
        RECT 0.1419 0.13 0.146 0.23 ;
        RECT 0.1419 0.23 0.146 0.25 ;
        RECT 0.1419 0.25 0.146 0.258 ;
        RECT 0.146 0.1019 0.17 0.13 ;
        RECT 0.146 0.13 0.17 0.23 ;
        RECT 0.146 0.23 0.17 0.25 ;
        RECT 0.146 0.25 0.17 0.258 ;
        RECT 0.146 0.574 0.17 0.602 ;
        RECT 0.17 0.1019 0.306 0.13 ;
        RECT 0.17 0.23 0.306 0.25 ;
        RECT 0.17 0.25 0.306 0.258 ;
        RECT 0.17 0.574 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.25 ;
        RECT 0.306 0.25 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.294 ;
        RECT 0.306 0.294 0.334 0.574 ;
        RECT 0.306 0.574 0.334 0.602 ;
        RECT 0.334 0.1019 0.782 0.13 ;
        RECT 0.782 0.1019 0.8139 0.13 ;
        RECT 0.782 0.13 0.8139 0.23 ;
        RECT 0.782 0.23 0.8139 0.25 ;
        RECT 0.782 0.25 0.8139 0.258 ;
        RECT 0.782 0.258 0.8139 0.294 ;
        RECT 0.8139 0.25 1.593 0.258 ;
        RECT 0.8139 0.258 1.593 0.294 ;
      LAYER M1 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.356 ;
        RECT 0.37 0.356 0.398 0.378 ;
        RECT 0.37 0.378 0.398 0.426 ;
        RECT 0.37 0.426 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.783 0.666 ;
        RECT 0.783 0.356 0.839 0.378 ;
        RECT 0.783 0.378 0.839 0.426 ;
        RECT 0.783 0.426 0.839 0.638 ;
        RECT 0.783 0.638 0.839 0.666 ;
        RECT 0.839 0.378 1.557 0.426 ;
        RECT 0.882 0.1019 0.931 0.13 ;
        RECT 0.931 0.1019 0.989 0.13 ;
        RECT 0.931 0.532 0.989 0.5639 ;
        RECT 0.931 0.5639 0.989 0.62 ;
        RECT 0.989 0.1019 1.572 0.13 ;
        RECT 0.989 0.532 1.572 0.5639 ;
        RECT 1.572 0.073 1.586 0.1019 ;
        RECT 1.572 0.1019 1.586 0.13 ;
        RECT 1.572 0.532 1.586 0.5639 ;
        RECT 1.586 0.073 1.614 0.1019 ;
        RECT 1.586 0.1019 1.614 0.13 ;
        RECT 1.586 0.532 1.614 0.5639 ;
        RECT 1.586 0.5639 1.614 0.62 ;
        RECT 1.586 0.62 1.614 0.624 ;
        RECT 1.614 0.073 1.6279 0.1019 ;
        RECT 1.614 0.1019 1.6279 0.13 ;
        RECT 1.614 0.532 1.6279 0.5639 ;
        RECT 1.6279 0.1019 1.629 0.13 ;
        RECT 1.6279 0.532 1.629 0.5639 ;
        RECT 1.629 0.1019 1.684 0.13 ;
        RECT 1.629 0.13 1.684 0.532 ;
        RECT 1.629 0.532 1.684 0.5639 ;
        RECT 0.05 0.1739 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.672 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.1419 0.1019 0.146 0.13 ;
        RECT 0.1419 0.13 0.146 0.23 ;
        RECT 0.1419 0.23 0.146 0.25 ;
        RECT 0.1419 0.25 0.146 0.258 ;
        RECT 0.146 0.1019 0.17 0.13 ;
        RECT 0.146 0.13 0.17 0.23 ;
        RECT 0.146 0.23 0.17 0.25 ;
        RECT 0.146 0.25 0.17 0.258 ;
        RECT 0.146 0.574 0.17 0.602 ;
        RECT 0.17 0.1019 0.306 0.13 ;
        RECT 0.17 0.23 0.306 0.25 ;
        RECT 0.17 0.25 0.306 0.258 ;
        RECT 0.17 0.574 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.25 ;
        RECT 0.306 0.25 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.294 ;
        RECT 0.306 0.294 0.334 0.574 ;
        RECT 0.306 0.574 0.334 0.602 ;
        RECT 0.334 0.1019 0.782 0.13 ;
        RECT 0.782 0.1019 0.8139 0.13 ;
        RECT 0.782 0.13 0.8139 0.23 ;
        RECT 0.782 0.23 0.8139 0.25 ;
        RECT 0.782 0.25 0.8139 0.258 ;
        RECT 0.782 0.258 0.8139 0.294 ;
        RECT 0.8139 0.25 1.593 0.258 ;
        RECT 0.8139 0.258 1.593 0.294 ;
  END
END TBUF_X12_12T

MACRO TBUF_X16_12T
  CLASS core ;
  FOREIGN TBUF_X16_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 3.168 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.39 0.1419 0.486 ;
        RECT 0.114 0.486 0.1419 0.514 ;
        RECT 0.1419 0.486 0.1739 0.514 ;
        RECT 0.1739 0.486 0.24 0.514 ;
        RECT 0.24 0.32 0.272 0.39 ;
        RECT 0.24 0.39 0.272 0.486 ;
        RECT 0.24 0.486 0.272 0.514 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.462 0.402 0.562 0.448 ;
        RECT 0.562 0.3459 0.59 0.402 ;
        RECT 0.562 0.402 0.59 0.448 ;
        RECT 0.59 0.402 0.6899 0.448 ;
        RECT 0.6899 0.402 0.718 0.448 ;
        RECT 0.6899 0.448 0.718 0.576 ;
        RECT 0.718 0.402 0.902 0.448 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.072 0.064 1.104 0.1419 ;
        RECT 1.072 0.1419 1.104 0.2 ;
        RECT 1.072 0.52 1.104 0.576 ;
        RECT 1.072 0.576 1.104 0.704 ;
        RECT 1.104 0.1419 1.968 0.2 ;
        RECT 1.104 0.52 1.968 0.576 ;
        RECT 1.968 0.064 1.98 0.1419 ;
        RECT 1.968 0.1419 1.98 0.2 ;
        RECT 1.968 0.52 1.98 0.576 ;
        RECT 1.968 0.576 1.98 0.704 ;
        RECT 1.98 0.064 1.998 0.1419 ;
        RECT 1.98 0.1419 1.998 0.2 ;
        RECT 1.98 0.52 1.998 0.576 ;
        RECT 1.98 0.576 1.998 0.704 ;
        RECT 1.998 0.064 2 0.1419 ;
        RECT 1.998 0.1419 2 0.2 ;
        RECT 1.998 0.52 2 0.576 ;
        RECT 1.998 0.576 2 0.704 ;
        RECT 2 0.1419 2.0339 0.2 ;
        RECT 2 0.52 2.0339 0.576 ;
        RECT 2.0339 0.1419 2.062 0.2 ;
        RECT 2.0339 0.2 2.062 0.52 ;
        RECT 2.0339 0.52 2.062 0.576 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.98 0.796 ;
        RECT 1.98 0.74 1.998 0.796 ;
        RECT 1.998 0.74 2.122 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 2.122 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.262 ;
        RECT 0.05 0.262 0.078 0.29 ;
        RECT 0.05 0.29 0.078 0.3459 ;
        RECT 0.05 0.3459 0.078 0.6 ;
        RECT 0.078 0.262 0.1419 0.29 ;
        RECT 0.1419 0.262 0.1739 0.29 ;
        RECT 0.1419 0.29 0.1739 0.3459 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.398 0.198 ;
        RECT 0.274 0.638 0.398 0.666 ;
        RECT 0.398 0.166 0.426 0.198 ;
        RECT 0.398 0.198 0.426 0.403 ;
        RECT 0.398 0.403 0.426 0.461 ;
        RECT 0.398 0.461 0.426 0.638 ;
        RECT 0.398 0.638 0.426 0.666 ;
        RECT 0.426 0.638 0.946 0.666 ;
        RECT 0.946 0.403 0.974 0.461 ;
        RECT 0.946 0.461 0.974 0.638 ;
        RECT 0.946 0.638 0.974 0.666 ;
        RECT 0.974 0.403 1.98 0.461 ;
        RECT 0.146 0.5679 0.21 0.602 ;
        RECT 0.21 0.1019 0.238 0.13 ;
        RECT 0.21 0.13 0.238 0.234 ;
        RECT 0.21 0.234 0.238 0.262 ;
        RECT 0.21 0.5679 0.238 0.602 ;
        RECT 0.238 0.1019 0.326 0.13 ;
        RECT 0.238 0.234 0.326 0.262 ;
        RECT 0.238 0.5679 0.326 0.602 ;
        RECT 0.326 0.1019 0.362 0.13 ;
        RECT 0.326 0.234 0.362 0.262 ;
        RECT 0.326 0.262 0.362 0.273 ;
        RECT 0.326 0.273 0.362 0.331 ;
        RECT 0.326 0.331 0.362 0.5679 ;
        RECT 0.326 0.5679 0.362 0.602 ;
        RECT 0.362 0.1019 0.946 0.13 ;
        RECT 0.946 0.1019 0.974 0.13 ;
        RECT 0.946 0.13 0.974 0.234 ;
        RECT 0.946 0.234 0.974 0.262 ;
        RECT 0.946 0.262 0.974 0.273 ;
        RECT 0.946 0.273 0.974 0.331 ;
        RECT 0.974 0.273 1.998 0.331 ;
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.262 ;
        RECT 0.05 0.262 0.078 0.29 ;
        RECT 0.05 0.29 0.078 0.3459 ;
        RECT 0.05 0.3459 0.078 0.6 ;
        RECT 0.078 0.262 0.1419 0.29 ;
        RECT 0.1419 0.262 0.1739 0.29 ;
        RECT 0.1419 0.29 0.1739 0.3459 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.398 0.198 ;
        RECT 0.274 0.638 0.398 0.666 ;
        RECT 0.398 0.166 0.426 0.198 ;
        RECT 0.398 0.198 0.426 0.403 ;
        RECT 0.398 0.403 0.426 0.461 ;
        RECT 0.398 0.461 0.426 0.638 ;
        RECT 0.398 0.638 0.426 0.666 ;
        RECT 0.426 0.638 0.946 0.666 ;
        RECT 0.946 0.403 0.974 0.461 ;
        RECT 0.946 0.461 0.974 0.638 ;
        RECT 0.946 0.638 0.974 0.666 ;
        RECT 0.974 0.403 1.98 0.461 ;
        RECT 0.146 0.5679 0.21 0.602 ;
        RECT 0.21 0.1019 0.238 0.13 ;
        RECT 0.21 0.13 0.238 0.234 ;
        RECT 0.21 0.234 0.238 0.262 ;
        RECT 0.21 0.5679 0.238 0.602 ;
        RECT 0.238 0.1019 0.326 0.13 ;
        RECT 0.238 0.234 0.326 0.262 ;
        RECT 0.238 0.5679 0.326 0.602 ;
        RECT 0.326 0.1019 0.362 0.13 ;
        RECT 0.326 0.234 0.362 0.262 ;
        RECT 0.326 0.262 0.362 0.273 ;
        RECT 0.326 0.273 0.362 0.331 ;
        RECT 0.326 0.331 0.362 0.5679 ;
        RECT 0.326 0.5679 0.362 0.602 ;
        RECT 0.362 0.1019 0.946 0.13 ;
        RECT 0.946 0.1019 0.974 0.13 ;
        RECT 0.946 0.13 0.974 0.234 ;
        RECT 0.946 0.234 0.974 0.262 ;
        RECT 0.946 0.262 0.974 0.273 ;
        RECT 0.946 0.273 0.974 0.331 ;
        RECT 0.974 0.273 1.998 0.331 ;
  END
END TBUF_X16_12T

MACRO TIEH_12T
  CLASS core ;
  FOREIGN TIEH_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.288 BY 0.512 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.473 0.1419 0.704 ;
        RECT 0.1419 0.473 0.147 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.096 0.1419 0.429 ;
      LAYER M1 ;
        RECT 0.114 0.096 0.1419 0.429 ;
  END
END TIEH_12T

MACRO TIEL_12T
  CLASS core ;
  FOREIGN TIEL_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.288 BY 0.512 ;
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.064 0.147 0.266 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.336 0.1419 0.672 ;
      LAYER M1 ;
        RECT 0.114 0.336 0.1419 0.672 ;
  END
END TIEL_12T

MACRO XNOR2_X1_12T
  CLASS core ;
  FOREIGN XNOR2_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.252 0.21 0.28 ;
        RECT 0.178 0.28 0.21 0.428 ;
        RECT 0.21 0.252 0.37 0.28 ;
        RECT 0.37 0.252 0.398 0.28 ;
        RECT 0.37 0.28 0.398 0.428 ;
        RECT 0.37 0.428 0.398 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.242 0.078 0.32 ;
        RECT 0.05 0.32 0.078 0.676 ;
        RECT 0.05 0.676 0.078 0.704 ;
        RECT 0.078 0.676 0.274 0.704 ;
        RECT 0.274 0.676 0.498 0.704 ;
        RECT 0.498 0.32 0.526 0.676 ;
        RECT 0.498 0.676 0.526 0.704 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.278 0.546 0.302 0.547 ;
        RECT 0.278 0.547 0.302 0.601 ;
        RECT 0.278 0.601 0.302 0.602 ;
        RECT 0.302 0.166 0.334 0.194 ;
        RECT 0.302 0.546 0.334 0.547 ;
        RECT 0.302 0.547 0.334 0.601 ;
        RECT 0.302 0.601 0.334 0.602 ;
        RECT 0.334 0.166 0.434 0.194 ;
        RECT 0.334 0.547 0.434 0.601 ;
        RECT 0.434 0.166 0.462 0.194 ;
        RECT 0.434 0.248 0.462 0.276 ;
        RECT 0.434 0.276 0.462 0.546 ;
        RECT 0.434 0.546 0.462 0.547 ;
        RECT 0.434 0.547 0.462 0.601 ;
        RECT 0.462 0.166 0.493 0.194 ;
        RECT 0.462 0.248 0.493 0.276 ;
        RECT 0.493 0.166 0.531 0.194 ;
        RECT 0.493 0.194 0.531 0.248 ;
        RECT 0.493 0.248 0.531 0.276 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.274 0.796 ;
        RECT 0.274 0.74 0.535 0.796 ;
        RECT 0.535 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.1019 0.535 0.13 ;
        RECT 0.114 0.184 0.1419 0.216 ;
        RECT 0.114 0.216 0.1419 0.34 ;
        RECT 0.114 0.34 0.1419 0.464 ;
        RECT 0.114 0.464 0.1419 0.492 ;
        RECT 0.114 0.492 0.1419 0.552 ;
        RECT 0.1419 0.184 0.234 0.216 ;
        RECT 0.1419 0.464 0.234 0.492 ;
        RECT 0.234 0.464 0.246 0.492 ;
        RECT 0.246 0.34 0.274 0.464 ;
        RECT 0.246 0.464 0.274 0.492 ;
      LAYER M1 ;
        RECT 0.21 0.1019 0.535 0.13 ;
        RECT 0.114 0.184 0.1419 0.216 ;
        RECT 0.114 0.216 0.1419 0.34 ;
        RECT 0.114 0.34 0.1419 0.464 ;
        RECT 0.114 0.464 0.1419 0.492 ;
        RECT 0.114 0.492 0.1419 0.552 ;
        RECT 0.1419 0.184 0.234 0.216 ;
        RECT 0.1419 0.464 0.234 0.492 ;
        RECT 0.234 0.464 0.246 0.492 ;
        RECT 0.246 0.34 0.274 0.464 ;
        RECT 0.246 0.464 0.274 0.492 ;
  END
END XNOR2_X1_12T

MACRO XOR2_X1_12T
  CLASS core ;
  FOREIGN XOR2_X1_12T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.864 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.3439 0.21 0.486 ;
        RECT 0.178 0.486 0.21 0.514 ;
        RECT 0.21 0.486 0.274 0.514 ;
        RECT 0.274 0.486 0.37 0.514 ;
        RECT 0.37 0.32 0.398 0.3439 ;
        RECT 0.37 0.3439 0.398 0.486 ;
        RECT 0.37 0.486 0.398 0.514 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.064 0.078 0.092 ;
        RECT 0.05 0.092 0.078 0.448 ;
        RECT 0.05 0.448 0.078 0.526 ;
        RECT 0.078 0.064 0.498 0.092 ;
        RECT 0.498 0.064 0.526 0.092 ;
        RECT 0.498 0.092 0.526 0.448 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.275 0.163 0.315 0.164 ;
        RECT 0.275 0.164 0.315 0.222 ;
        RECT 0.315 0.163 0.334 0.164 ;
        RECT 0.315 0.164 0.334 0.222 ;
        RECT 0.315 0.574 0.334 0.602 ;
        RECT 0.334 0.164 0.434 0.222 ;
        RECT 0.334 0.574 0.434 0.602 ;
        RECT 0.434 0.164 0.462 0.222 ;
        RECT 0.434 0.222 0.462 0.492 ;
        RECT 0.434 0.492 0.462 0.52 ;
        RECT 0.434 0.574 0.462 0.602 ;
        RECT 0.462 0.492 0.496 0.52 ;
        RECT 0.462 0.574 0.496 0.602 ;
        RECT 0.496 0.492 0.528 0.52 ;
        RECT 0.496 0.52 0.528 0.574 ;
        RECT 0.496 0.574 0.528 0.602 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.535 0.796 ;
        RECT 0.535 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.246 0.638 0.535 0.666 ;
        RECT 0.114 0.136 0.1419 0.28 ;
        RECT 0.114 0.28 0.1419 0.308 ;
        RECT 0.114 0.308 0.1419 0.432 ;
        RECT 0.114 0.432 0.1419 0.552 ;
        RECT 0.114 0.552 0.1419 0.584 ;
        RECT 0.1419 0.28 0.246 0.308 ;
        RECT 0.1419 0.552 0.246 0.584 ;
        RECT 0.246 0.28 0.247 0.308 ;
        RECT 0.246 0.308 0.247 0.432 ;
        RECT 0.246 0.552 0.247 0.584 ;
        RECT 0.247 0.28 0.274 0.308 ;
        RECT 0.247 0.308 0.274 0.432 ;
      LAYER M1 ;
        RECT 0.246 0.638 0.535 0.666 ;
        RECT 0.114 0.136 0.1419 0.28 ;
        RECT 0.114 0.28 0.1419 0.308 ;
        RECT 0.114 0.308 0.1419 0.432 ;
        RECT 0.114 0.432 0.1419 0.552 ;
        RECT 0.114 0.552 0.1419 0.584 ;
        RECT 0.1419 0.28 0.246 0.308 ;
        RECT 0.1419 0.552 0.246 0.584 ;
        RECT 0.246 0.28 0.247 0.308 ;
        RECT 0.246 0.308 0.247 0.432 ;
        RECT 0.246 0.552 0.247 0.584 ;
        RECT 0.247 0.28 0.274 0.308 ;
        RECT 0.247 0.308 0.274 0.432 ;
  END
END XOR2_X1_12T

END LIBRARY
#
# End of file
#
